`timescale 1ns/1ps
module tb;
    localparam int N_INPUTS = 10;
    localparam int OUT_WIDTH = 11;
    localparam logic [(11264)-1:0] TT = 11264'h5A4B4D49E935A4B4D69A935A4B6D6DADB1B4B6D6DAFB584B4F49E93584B4D69E931A4B4D69ADB1B436C6DAFBD85B0F41E93184B0F69E9318430C69EF318434C7D8FB985B0F41E8798530E61E8318430E61CF338430C71CF3584B4949A93584B4969A935A4B4969ADB1B43696DAFB584B0941E93584B0969A9318430969AF31843487DAFB585B0B41E8718430961E8318430861AF3384308718F398530B43E8718530A61EA738430871CE7384788718E7584B0941292584B0969292184B09692F23843497D2FA584B0941286184B0961282184309612F2384708710F2184B0B43686184309612A6384308710E6384788F10E618531B4368638430A634A6384708730E6384788F31E6584B0941286584B0961282384B09612F2384708712F2584B0943286184B09612A6384708712E6384788F10E6184B1943686384308632A6384708F30E6384788F31E638C31A436A6384718734A6384798F31E63C4798F31E65A6B4F49E935A6B4D6DA9B5B6B6D6DA9B5B6B6D6DADB5A7B4F49E935A6B4F69E935A6B6D6DA9B1B636D6DADBD87B0F49E93587B4F69E9318634F69E9B1B636C6DAFBD87B0F41E9398730F61E9318730E69E9318630E6DCFB5A4B4D49E935A4B4D69A935A4B6D6DA9B1B4B6D6DADB584B0F49E93584B4D69E93184B4D69A9B1B436D6DAFBD85B0F41E93184B0F61E9318430D69E9338430C6D8FB985B0F41E8798530F61E8718430E61CA338470C71CF3584B0949293584B4969293584B496929B1B4B696D2FB584B0941693584B0961293184B09692933843086D2FB585B0B41687184B0961687384308612A3384708710F3985B0B4368718530A63687384708614A7384708F10E7584B0941292584B0961292584B09692923847096D2FA584B0941286584B0961286384309612A2384708F12F2584B0B4368638430963286384708612A6384708F11E618531B4368638471A636A6384708F30A6384788F31E65A7B4F49E9B5B6B6D4DE9B5B6B6D6DA9B5B6B6D6DA5BDA7B4F49E935A7B4F4DE9B5B6B6D6DE9B1B6B6D6DA5BD87B4F49E93DA7B4F49E931A7B6F6DE9B1B636D6DE5BD87B0F49E93987B0F49E9398734F69E9B19736E6DC5B5A6B4F49E935A6B4D4DA9B5B6B6D6DA9B5B6B6D6DADB587B4F49E935A6B4F49E935A6B6D6DA9B1B6B6D6DADBD87B0F49E93587B0F49E93186B4F69E9B19636C6DADBD87B0F41E83987B0F41E9318730E61E9338630E6DCFB584B4949E935A4B4949A935A4B696DA9B5B4B696DADB584B0B49E93584B0949E93584B4969A9B3943696DADBD85B0B41E83584B0B41E9318430961E933847086DAFBD85B0B41E8798530B41E8738430A61E87384708E1CE3584B0949293584B0949293584B496929B394B696D2DB584B0941683584B0941293384B09612933847096D2FB585B0B41687184B094168738470961287384708E10E3985B0B4368738530B43687384708E34A7384708F11E7DA7A6F4DE9B5B6B6F4DE9B5B6B6D6DE1B5B6B6D2DA1BDA7A4F49E9BDB7B6F4DE9B5B6B6F6DE1B5B6B6D2DE1BDA7A4F49E93DA7B4F4DE9BDB7B6F6DE1B1B6B6F2DE1BD87A4F49E93D87B4F49E939A7B6F6DE1B9B736E2DE1B5A7A4F49E9B5B6B6D4DE9B5B6B6D6DA9B5B6B6D6DA1BDA7A4F49E935A7B4F4DE9B5B6B6D6DE9B5B6B6D6DA1BD87A4F49E93D87B4F49E935A7B6F6DE9B1B636D6DE1BD87A0F41E93D87B0F49E9398730F69E9B39736E6DE1B5A4A4F49E935A4B4D4DA9B5B4B6D6DA9B5B4B6D6DA9B585A4F49E93584B4F49E935A4B6D6DA9B1B4B6D6DA9BD85A0F41E93585B0F49E93184B0F69E9B39436D6DA9BD85A0F41E87985B0F41E8338530F61E9338470E65C9B584A4949E93584B4949A935A4B696DA9B7B4B696DA9B584A0B41E93584B0949E93584B0969A9B394F696DA9BD85A0B41E87584B0B41E83384B0961E93384708E5A9BD85A0B43E87B85B0B41E8738470A61E87384708E1DA7;
    reg  [N_INPUTS-1:0] x;
    wire [OUT_WIDTH-1:0] f;

    top dut (.x(x), .f(f));

    integer i;
    initial begin
        for (i = 0; i < (1<<N_INPUTS); i = i + 1) begin
            x = i[N_INPUTS-1:0];
            #1;
            if (f !== TT[i*OUT_WIDTH +: OUT_WIDTH]) begin
                $error("Mismatch at %0d: expected %0b got %0b", i, TT[i*OUT_WIDTH +: OUT_WIDTH], f);
                $finish;
            end
        end
        $display("PASS: all patterns matched.");
        $finish;
    end
endmodule
