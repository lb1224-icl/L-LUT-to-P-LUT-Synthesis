`timescale 1ns/1ps
module top (input wire [11:0] x, output wire [11:0] f);
    (* KEEP = "TRUE" *) wire n0;
    (* KEEP = "TRUE" *) wire n1;
    (* KEEP = "TRUE" *) wire n2;
    (* KEEP = "TRUE" *) wire n3;
    (* KEEP = "TRUE" *) wire n4;
    (* KEEP = "TRUE" *) wire n5;
    (* KEEP = "TRUE" *) wire n6;
    (* KEEP = "TRUE" *) wire n7;
    (* KEEP = "TRUE" *) wire n8;
    (* KEEP = "TRUE" *) wire n9;
    (* KEEP = "TRUE" *) wire n10;
    (* KEEP = "TRUE" *) wire n11;
    (* KEEP = "TRUE" *) wire n12;
    (* KEEP = "TRUE" *) wire n13;
    (* KEEP = "TRUE" *) wire n14;
    (* KEEP = "TRUE" *) wire n15;
    (* KEEP = "TRUE" *) wire n16;
    (* KEEP = "TRUE" *) wire n17;
    (* KEEP = "TRUE" *) wire n18;
    (* KEEP = "TRUE" *) wire n19;
    (* KEEP = "TRUE" *) wire n20;
    (* KEEP = "TRUE" *) wire n21;
    (* KEEP = "TRUE" *) wire n22;
    (* KEEP = "TRUE" *) wire n23;
    (* KEEP = "TRUE" *) wire n24;
    (* KEEP = "TRUE" *) wire n25;
    (* KEEP = "TRUE" *) wire n26;
    (* KEEP = "TRUE" *) wire n27;
    (* KEEP = "TRUE" *) wire n28;
    (* KEEP = "TRUE" *) wire n29;
    (* KEEP = "TRUE" *) wire n30;
    (* KEEP = "TRUE" *) wire n31;
    (* KEEP = "TRUE" *) wire n32;
    (* KEEP = "TRUE" *) wire n33;
    (* KEEP = "TRUE" *) wire n34;
    (* KEEP = "TRUE" *) wire n35;
    (* KEEP = "TRUE" *) wire n36;
    (* KEEP = "TRUE" *) wire n37;
    (* KEEP = "TRUE" *) wire n38;
    (* KEEP = "TRUE" *) wire n39;
    (* KEEP = "TRUE" *) wire n40;
    (* KEEP = "TRUE" *) wire n41;
    (* KEEP = "TRUE" *) wire n42;
    (* KEEP = "TRUE" *) wire n43;
    (* KEEP = "TRUE" *) wire n44;
    (* KEEP = "TRUE" *) wire n45;
    (* KEEP = "TRUE" *) wire n46;
    (* KEEP = "TRUE" *) wire n47;
    (* KEEP = "TRUE" *) wire n48;
    (* KEEP = "TRUE" *) wire n49;
    (* KEEP = "TRUE" *) wire n50;
    (* KEEP = "TRUE" *) wire n51;
    (* KEEP = "TRUE" *) wire n52;
    (* KEEP = "TRUE" *) wire n53;
    (* KEEP = "TRUE" *) wire n54;
    (* KEEP = "TRUE" *) wire n55;
    (* KEEP = "TRUE" *) wire n56;
    (* KEEP = "TRUE" *) wire n57;
    (* KEEP = "TRUE" *) wire n58;
    (* KEEP = "TRUE" *) wire n59;
    (* KEEP = "TRUE" *) wire n60;
    (* KEEP = "TRUE" *) wire n61;
    (* KEEP = "TRUE" *) wire n62;
    (* KEEP = "TRUE" *) wire n63;
    (* KEEP = "TRUE" *) wire n64;
    (* KEEP = "TRUE" *) wire n65;
    (* KEEP = "TRUE" *) wire n66;
    (* KEEP = "TRUE" *) wire n67;
    (* KEEP = "TRUE" *) wire n68;
    (* KEEP = "TRUE" *) wire n69;
    (* KEEP = "TRUE" *) wire n70;
    (* KEEP = "TRUE" *) wire n71;
    (* KEEP = "TRUE" *) wire n72;
    (* KEEP = "TRUE" *) wire n73;
    (* KEEP = "TRUE" *) wire n74;
    (* KEEP = "TRUE" *) wire n75;
    (* KEEP = "TRUE" *) wire n76;
    (* KEEP = "TRUE" *) wire n77;
    (* KEEP = "TRUE" *) wire n78;
    (* KEEP = "TRUE" *) wire n79;
    (* KEEP = "TRUE" *) wire n80;
    (* KEEP = "TRUE" *) wire n81;
    (* KEEP = "TRUE" *) wire n82;
    (* KEEP = "TRUE" *) wire n83;
    (* KEEP = "TRUE" *) wire n84;
    (* KEEP = "TRUE" *) wire n85;
    (* KEEP = "TRUE" *) wire n86;
    (* KEEP = "TRUE" *) wire n87;
    (* KEEP = "TRUE" *) wire n88;
    (* KEEP = "TRUE" *) wire n89;
    (* KEEP = "TRUE" *) wire n90;
    (* KEEP = "TRUE" *) wire n91;
    (* KEEP = "TRUE" *) wire n92;
    (* KEEP = "TRUE" *) wire n93;
    (* KEEP = "TRUE" *) wire n94;
    (* KEEP = "TRUE" *) wire n95;
    (* KEEP = "TRUE" *) wire n96;
    (* KEEP = "TRUE" *) wire n97;
    (* KEEP = "TRUE" *) wire n98;
    (* KEEP = "TRUE" *) wire n99;
    (* KEEP = "TRUE" *) wire n100;
    (* KEEP = "TRUE" *) wire n101;
    (* KEEP = "TRUE" *) wire n102;
    (* KEEP = "TRUE" *) wire n103;
    (* KEEP = "TRUE" *) wire n104;
    (* KEEP = "TRUE" *) wire n105;
    (* KEEP = "TRUE" *) wire n106;
    (* KEEP = "TRUE" *) wire n107;
    (* KEEP = "TRUE" *) wire n108;
    (* KEEP = "TRUE" *) wire n109;
    (* KEEP = "TRUE" *) wire n110;
    (* KEEP = "TRUE" *) wire n111;
    (* KEEP = "TRUE" *) wire n112;
    (* KEEP = "TRUE" *) wire n113;
    (* KEEP = "TRUE" *) wire n114;
    (* KEEP = "TRUE" *) wire n115;
    (* KEEP = "TRUE" *) wire n116;
    (* KEEP = "TRUE" *) wire n117;
    (* KEEP = "TRUE" *) wire n118;
    (* KEEP = "TRUE" *) wire n119;
    (* KEEP = "TRUE" *) wire n120;
    (* KEEP = "TRUE" *) wire n121;
    (* KEEP = "TRUE" *) wire n122;
    (* KEEP = "TRUE" *) wire n123;
    (* KEEP = "TRUE" *) wire n124;
    (* KEEP = "TRUE" *) wire n125;
    (* KEEP = "TRUE" *) wire n126;
    (* KEEP = "TRUE" *) wire n127;
    (* KEEP = "TRUE" *) wire n128;
    (* KEEP = "TRUE" *) wire n129;
    (* KEEP = "TRUE" *) wire n130;
    (* KEEP = "TRUE" *) wire n131;
    (* KEEP = "TRUE" *) wire n132;
    (* KEEP = "TRUE" *) wire n133;
    (* KEEP = "TRUE" *) wire n134;
    (* KEEP = "TRUE" *) wire n135;
    (* KEEP = "TRUE" *) wire n136;
    (* KEEP = "TRUE" *) wire n137;
    (* KEEP = "TRUE" *) wire n138;
    (* KEEP = "TRUE" *) wire n139;
    (* KEEP = "TRUE" *) wire n140;
    (* KEEP = "TRUE" *) wire n141;
    (* KEEP = "TRUE" *) wire n142;
    (* KEEP = "TRUE" *) wire n143;
    (* KEEP = "TRUE" *) wire n144;
    (* KEEP = "TRUE" *) wire n145;
    (* KEEP = "TRUE" *) wire n146;
    (* KEEP = "TRUE" *) wire n147;
    (* KEEP = "TRUE" *) wire n148;
    (* KEEP = "TRUE" *) wire n149;
    (* KEEP = "TRUE" *) wire n150;
    (* KEEP = "TRUE" *) wire n151;
    (* KEEP = "TRUE" *) wire n152;
    (* KEEP = "TRUE" *) wire n153;
    (* KEEP = "TRUE" *) wire n154;
    (* KEEP = "TRUE" *) wire n155;
    (* KEEP = "TRUE" *) wire n156;
    (* KEEP = "TRUE" *) wire n157;
    (* KEEP = "TRUE" *) wire n158;
    (* KEEP = "TRUE" *) wire n159;
    (* KEEP = "TRUE" *) wire n160;
    (* KEEP = "TRUE" *) wire n161;
    (* KEEP = "TRUE" *) wire n162;
    (* KEEP = "TRUE" *) wire n163;
    (* KEEP = "TRUE" *) wire n164;
    (* KEEP = "TRUE" *) wire n165;
    (* KEEP = "TRUE" *) wire n166;
    (* KEEP = "TRUE" *) wire n167;
    (* KEEP = "TRUE" *) wire n168;
    (* KEEP = "TRUE" *) wire n169;
    (* KEEP = "TRUE" *) wire n170;
    (* KEEP = "TRUE" *) wire n171;
    (* KEEP = "TRUE" *) wire n172;
    (* KEEP = "TRUE" *) wire n173;
    (* KEEP = "TRUE" *) wire n174;
    (* KEEP = "TRUE" *) wire n175;
    (* KEEP = "TRUE" *) wire n176;
    (* KEEP = "TRUE" *) wire n177;
    (* KEEP = "TRUE" *) wire n178;
    (* KEEP = "TRUE" *) wire n179;
    (* KEEP = "TRUE" *) wire n180;
    (* KEEP = "TRUE" *) wire n181;
    (* KEEP = "TRUE" *) wire n182;
    (* KEEP = "TRUE" *) wire n183;
    (* KEEP = "TRUE" *) wire n184;
    (* KEEP = "TRUE" *) wire n185;
    (* KEEP = "TRUE" *) wire n186;
    (* KEEP = "TRUE" *) wire n187;
    (* KEEP = "TRUE" *) wire n188;
    (* KEEP = "TRUE" *) wire n189;
    (* KEEP = "TRUE" *) wire n190;
    (* KEEP = "TRUE" *) wire n191;
    (* KEEP = "TRUE" *) wire n192;
    (* KEEP = "TRUE" *) wire n193;
    (* KEEP = "TRUE" *) wire n194;
    (* KEEP = "TRUE" *) wire n195;
    (* KEEP = "TRUE" *) wire n196;
    (* KEEP = "TRUE" *) wire n197;
    (* KEEP = "TRUE" *) wire n198;
    (* KEEP = "TRUE" *) wire n199;
    (* KEEP = "TRUE" *) wire n200;
    (* KEEP = "TRUE" *) wire n201;
    (* KEEP = "TRUE" *) wire n202;
    (* KEEP = "TRUE" *) wire n203;
    (* KEEP = "TRUE" *) wire n204;
    (* KEEP = "TRUE" *) wire n205;
    (* KEEP = "TRUE" *) wire n206;
    (* KEEP = "TRUE" *) wire n207;
    (* KEEP = "TRUE" *) wire n208;
    (* KEEP = "TRUE" *) wire n209;
    (* KEEP = "TRUE" *) wire n210;
    (* KEEP = "TRUE" *) wire n211;
    (* KEEP = "TRUE" *) wire n212;
    (* KEEP = "TRUE" *) wire n213;
    (* KEEP = "TRUE" *) wire n214;
    (* KEEP = "TRUE" *) wire n215;
    (* KEEP = "TRUE" *) wire n216;
    (* KEEP = "TRUE" *) wire n217;
    (* KEEP = "TRUE" *) wire n218;
    (* KEEP = "TRUE" *) wire n219;
    (* KEEP = "TRUE" *) wire n220;
    (* KEEP = "TRUE" *) wire n221;
    (* KEEP = "TRUE" *) wire n222;
    (* KEEP = "TRUE" *) wire n223;
    (* KEEP = "TRUE" *) wire n224;
    (* KEEP = "TRUE" *) wire n225;
    (* KEEP = "TRUE" *) wire n226;
    (* KEEP = "TRUE" *) wire n227;
    (* KEEP = "TRUE" *) wire n228;
    (* KEEP = "TRUE" *) wire n229;
    (* KEEP = "TRUE" *) wire n230;
    (* KEEP = "TRUE" *) wire n231;
    (* KEEP = "TRUE" *) wire n232;
    (* KEEP = "TRUE" *) wire n233;
    (* KEEP = "TRUE" *) wire n234;
    (* KEEP = "TRUE" *) wire n235;
    (* KEEP = "TRUE" *) wire n236;
    (* KEEP = "TRUE" *) wire n237;
    (* KEEP = "TRUE" *) wire n238;
    (* KEEP = "TRUE" *) wire n239;
    (* KEEP = "TRUE" *) wire n240;
    (* KEEP = "TRUE" *) wire n241;
    (* KEEP = "TRUE" *) wire n242;
    (* KEEP = "TRUE" *) wire n243;
    (* KEEP = "TRUE" *) wire n244;
    (* KEEP = "TRUE" *) wire n245;
    (* KEEP = "TRUE" *) wire n246;
    (* KEEP = "TRUE" *) wire n247;
    (* KEEP = "TRUE" *) wire n248;
    (* KEEP = "TRUE" *) wire n249;
    (* KEEP = "TRUE" *) wire n250;
    (* KEEP = "TRUE" *) wire n251;
    (* KEEP = "TRUE" *) wire n252;
    (* KEEP = "TRUE" *) wire n253;
    (* KEEP = "TRUE" *) wire n254;
    (* KEEP = "TRUE" *) wire n255;
    (* KEEP = "TRUE" *) wire n256;
    (* KEEP = "TRUE" *) wire n257;
    (* KEEP = "TRUE" *) wire n258;
    (* KEEP = "TRUE" *) wire n259;
    (* KEEP = "TRUE" *) wire n260;
    (* KEEP = "TRUE" *) wire n261;
    (* KEEP = "TRUE" *) wire n262;
    (* KEEP = "TRUE" *) wire n263;
    (* KEEP = "TRUE" *) wire n264;
    (* KEEP = "TRUE" *) wire n265;
    (* KEEP = "TRUE" *) wire n266;
    (* KEEP = "TRUE" *) wire n267;
    (* KEEP = "TRUE" *) wire n268;
    (* KEEP = "TRUE" *) wire n269;
    (* KEEP = "TRUE" *) wire n270;
    (* KEEP = "TRUE" *) wire n271;
    (* KEEP = "TRUE" *) wire n272;
    (* KEEP = "TRUE" *) wire n273;
    (* KEEP = "TRUE" *) wire n274;
    (* KEEP = "TRUE" *) wire n275;
    (* KEEP = "TRUE" *) wire n276;
    (* KEEP = "TRUE" *) wire n277;
    (* KEEP = "TRUE" *) wire n278;
    (* KEEP = "TRUE" *) wire n279;
    (* KEEP = "TRUE" *) wire n280;
    (* KEEP = "TRUE" *) wire n281;
    (* KEEP = "TRUE" *) wire n282;
    (* KEEP = "TRUE" *) wire n283;
    (* KEEP = "TRUE" *) wire n284;
    (* KEEP = "TRUE" *) wire n285;
    (* KEEP = "TRUE" *) wire n286;
    (* KEEP = "TRUE" *) wire n287;
    (* KEEP = "TRUE" *) wire n288;
    (* KEEP = "TRUE" *) wire n289;
    (* KEEP = "TRUE" *) wire n290;
    (* KEEP = "TRUE" *) wire n291;
    (* KEEP = "TRUE" *) wire n292;
    (* KEEP = "TRUE" *) wire n293;
    (* KEEP = "TRUE" *) wire n294;
    (* KEEP = "TRUE" *) wire n295;
    (* KEEP = "TRUE" *) wire n296;
    (* KEEP = "TRUE" *) wire n297;
    (* KEEP = "TRUE" *) wire n298;
    (* KEEP = "TRUE" *) wire n299;
    (* KEEP = "TRUE" *) wire n300;
    (* KEEP = "TRUE" *) wire n301;
    (* KEEP = "TRUE" *) wire n302;
    (* KEEP = "TRUE" *) wire n303;
    (* KEEP = "TRUE" *) wire n304;
    (* KEEP = "TRUE" *) wire n305;
    (* KEEP = "TRUE" *) wire n306;
    (* KEEP = "TRUE" *) wire n307;
    (* KEEP = "TRUE" *) wire n308;
    (* KEEP = "TRUE" *) wire n309;
    (* KEEP = "TRUE" *) wire n310;
    (* KEEP = "TRUE" *) wire n311;
    (* KEEP = "TRUE" *) wire n312;
    (* KEEP = "TRUE" *) wire n313;
    (* KEEP = "TRUE" *) wire n314;
    (* KEEP = "TRUE" *) wire n315;
    (* KEEP = "TRUE" *) wire n316;
    (* KEEP = "TRUE" *) wire n317;
    (* KEEP = "TRUE" *) wire n318;
    (* KEEP = "TRUE" *) wire n319;
    (* KEEP = "TRUE" *) wire n320;
    (* KEEP = "TRUE" *) wire n321;
    (* KEEP = "TRUE" *) wire n322;
    (* KEEP = "TRUE" *) wire n323;
    (* KEEP = "TRUE" *) wire n324;
    (* KEEP = "TRUE" *) wire n325;
    (* KEEP = "TRUE" *) wire n326;
    (* KEEP = "TRUE" *) wire n327;
    (* KEEP = "TRUE" *) wire n328;
    (* KEEP = "TRUE" *) wire n329;
    (* KEEP = "TRUE" *) wire n330;
    (* KEEP = "TRUE" *) wire n331;
    (* KEEP = "TRUE" *) wire n332;
    (* KEEP = "TRUE" *) wire n333;
    (* KEEP = "TRUE" *) wire n334;
    (* KEEP = "TRUE" *) wire n335;
    (* KEEP = "TRUE" *) wire n336;
    (* KEEP = "TRUE" *) wire n337;
    (* KEEP = "TRUE" *) wire n338;
    (* KEEP = "TRUE" *) wire n339;
    (* KEEP = "TRUE" *) wire n340;
    (* KEEP = "TRUE" *) wire n341;
    (* KEEP = "TRUE" *) wire n342;
    (* KEEP = "TRUE" *) wire n343;
    (* KEEP = "TRUE" *) wire n344;
    (* KEEP = "TRUE" *) wire n345;
    (* KEEP = "TRUE" *) wire n346;
    (* KEEP = "TRUE" *) wire n347;
    (* KEEP = "TRUE" *) wire n348;
    (* KEEP = "TRUE" *) wire n349;
    (* KEEP = "TRUE" *) wire n350;
    (* KEEP = "TRUE" *) wire n351;
    (* KEEP = "TRUE" *) wire n352;
    (* KEEP = "TRUE" *) wire n353;
    (* KEEP = "TRUE" *) wire n354;
    (* KEEP = "TRUE" *) wire n355;
    (* KEEP = "TRUE" *) wire n356;
    (* KEEP = "TRUE" *) wire n357;
    (* KEEP = "TRUE" *) wire n358;
    (* KEEP = "TRUE" *) wire n359;
    (* KEEP = "TRUE" *) wire n360;
    (* KEEP = "TRUE" *) wire n361;
    (* KEEP = "TRUE" *) wire n362;
    (* KEEP = "TRUE" *) wire n363;
    (* KEEP = "TRUE" *) wire n364;
    (* KEEP = "TRUE" *) wire n365;
    (* KEEP = "TRUE" *) wire n366;
    (* KEEP = "TRUE" *) wire n367;
    (* KEEP = "TRUE" *) wire n368;
    (* KEEP = "TRUE" *) wire n369;
    (* KEEP = "TRUE" *) wire n370;
    (* KEEP = "TRUE" *) wire n371;
    (* KEEP = "TRUE" *) wire n372;
    (* KEEP = "TRUE" *) wire n373;
    (* KEEP = "TRUE" *) wire n374;
    (* KEEP = "TRUE" *) wire n375;
    (* KEEP = "TRUE" *) wire n376;
    (* KEEP = "TRUE" *) wire n377;
    (* KEEP = "TRUE" *) wire n378;
    (* KEEP = "TRUE" *) wire n379;
    (* KEEP = "TRUE" *) wire n380;
    (* KEEP = "TRUE" *) wire n381;
    (* KEEP = "TRUE" *) wire n382;
    (* KEEP = "TRUE" *) wire n383;
    (* KEEP = "TRUE" *) wire n384;
    (* KEEP = "TRUE" *) wire n385;
    (* KEEP = "TRUE" *) wire n386;
    (* KEEP = "TRUE" *) wire n387;
    (* KEEP = "TRUE" *) wire n388;
    (* KEEP = "TRUE" *) wire n389;
    (* KEEP = "TRUE" *) wire n390;
    (* KEEP = "TRUE" *) wire n391;
    (* KEEP = "TRUE" *) wire n392;
    (* KEEP = "TRUE" *) wire n393;
    (* KEEP = "TRUE" *) wire n394;
    (* KEEP = "TRUE" *) wire n395;
    (* KEEP = "TRUE" *) wire n396;
    (* KEEP = "TRUE" *) wire n397;
    (* KEEP = "TRUE" *) wire n398;
    (* KEEP = "TRUE" *) wire n399;
    (* KEEP = "TRUE" *) wire n400;
    (* KEEP = "TRUE" *) wire n401;
    (* KEEP = "TRUE" *) wire n402;
    (* KEEP = "TRUE" *) wire n403;
    (* KEEP = "TRUE" *) wire n404;
    (* KEEP = "TRUE" *) wire n405;
    (* KEEP = "TRUE" *) wire n406;
    (* KEEP = "TRUE" *) wire n407;
    (* KEEP = "TRUE" *) wire n408;
    (* KEEP = "TRUE" *) wire n409;
    (* KEEP = "TRUE" *) wire n410;
    (* KEEP = "TRUE" *) wire n411;
    (* KEEP = "TRUE" *) wire n412;
    (* KEEP = "TRUE" *) wire n413;
    (* KEEP = "TRUE" *) wire n414;
    (* KEEP = "TRUE" *) wire n415;
    (* KEEP = "TRUE" *) wire n416;
    (* KEEP = "TRUE" *) wire n417;
    (* KEEP = "TRUE" *) wire n418;
    (* KEEP = "TRUE" *) wire n419;
    (* KEEP = "TRUE" *) wire n420;
    (* KEEP = "TRUE" *) wire n421;
    (* KEEP = "TRUE" *) wire n422;
    (* KEEP = "TRUE" *) wire n423;
    (* KEEP = "TRUE" *) wire n424;
    (* KEEP = "TRUE" *) wire n425;
    (* KEEP = "TRUE" *) wire n426;
    (* KEEP = "TRUE" *) wire n427;
    (* KEEP = "TRUE" *) wire n428;
    (* KEEP = "TRUE" *) wire n429;
    (* KEEP = "TRUE" *) wire n430;
    (* KEEP = "TRUE" *) wire n431;
    (* KEEP = "TRUE" *) wire n432;
    (* KEEP = "TRUE" *) wire n433;
    (* KEEP = "TRUE" *) wire n434;
    (* KEEP = "TRUE" *) wire n435;
    (* KEEP = "TRUE" *) wire n436;
    (* KEEP = "TRUE" *) wire n437;
    (* KEEP = "TRUE" *) wire n438;
    (* KEEP = "TRUE" *) wire n439;
    (* KEEP = "TRUE" *) wire n440;
    (* KEEP = "TRUE" *) wire n441;
    (* KEEP = "TRUE" *) wire n442;
    (* KEEP = "TRUE" *) wire n443;
    (* KEEP = "TRUE" *) wire n444;
    (* KEEP = "TRUE" *) wire n445;
    (* KEEP = "TRUE" *) wire n446;
    (* KEEP = "TRUE" *) wire n447;
    (* KEEP = "TRUE" *) wire n448;
    (* KEEP = "TRUE" *) wire n449;
    (* KEEP = "TRUE" *) wire n450;
    (* KEEP = "TRUE" *) wire n451;
    (* KEEP = "TRUE" *) wire n452;
    (* KEEP = "TRUE" *) wire n453;
    (* KEEP = "TRUE" *) wire n454;
    (* KEEP = "TRUE" *) wire n455;
    (* KEEP = "TRUE" *) wire n456;
    (* KEEP = "TRUE" *) wire n457;
    (* KEEP = "TRUE" *) wire n458;
    (* KEEP = "TRUE" *) wire n459;
    (* KEEP = "TRUE" *) wire n460;
    (* KEEP = "TRUE" *) wire n461;
    (* KEEP = "TRUE" *) wire n462;
    (* KEEP = "TRUE" *) wire n463;
    (* KEEP = "TRUE" *) wire n464;
    (* KEEP = "TRUE" *) wire n465;
    (* KEEP = "TRUE" *) wire n466;
    (* KEEP = "TRUE" *) wire n467;
    (* KEEP = "TRUE" *) wire n468;
    (* KEEP = "TRUE" *) wire n469;
    (* KEEP = "TRUE" *) wire n470;
    (* KEEP = "TRUE" *) wire n471;
    (* KEEP = "TRUE" *) wire n472;
    (* KEEP = "TRUE" *) wire n473;
    (* KEEP = "TRUE" *) wire n474;
    (* KEEP = "TRUE" *) wire n475;
    (* KEEP = "TRUE" *) wire n476;
    (* KEEP = "TRUE" *) wire n477;
    (* KEEP = "TRUE" *) wire n478;
    (* KEEP = "TRUE" *) wire n479;
    (* KEEP = "TRUE" *) wire n480;
    (* KEEP = "TRUE" *) wire n481;
    (* KEEP = "TRUE" *) wire n482;
    (* KEEP = "TRUE" *) wire n483;
    (* KEEP = "TRUE" *) wire n484;
    (* KEEP = "TRUE" *) wire n485;
    (* KEEP = "TRUE" *) wire n486;
    (* KEEP = "TRUE" *) wire n487;
    (* KEEP = "TRUE" *) wire n488;
    (* KEEP = "TRUE" *) wire n489;
    (* KEEP = "TRUE" *) wire n490;
    (* KEEP = "TRUE" *) wire n491;
    (* KEEP = "TRUE" *) wire n492;
    (* KEEP = "TRUE" *) wire n493;
    (* KEEP = "TRUE" *) wire n494;
    (* KEEP = "TRUE" *) wire n495;
    (* KEEP = "TRUE" *) wire n496;
    (* KEEP = "TRUE" *) wire n497;
    (* KEEP = "TRUE" *) wire n498;
    (* KEEP = "TRUE" *) wire n499;
    (* KEEP = "TRUE" *) wire n500;
    (* KEEP = "TRUE" *) wire n501;
    (* KEEP = "TRUE" *) wire n502;
    (* KEEP = "TRUE" *) wire n503;
    (* KEEP = "TRUE" *) wire n504;
    (* KEEP = "TRUE" *) wire n505;
    (* KEEP = "TRUE" *) wire n506;
    (* KEEP = "TRUE" *) wire n507;
    (* KEEP = "TRUE" *) wire n508;
    (* KEEP = "TRUE" *) wire n509;
    (* KEEP = "TRUE" *) wire n510;
    (* KEEP = "TRUE" *) wire n511;
    (* KEEP = "TRUE" *) wire n512;
    (* KEEP = "TRUE" *) wire n513;
    (* KEEP = "TRUE" *) wire n514;
    (* KEEP = "TRUE" *) wire n515;
    (* KEEP = "TRUE" *) wire n516;
    (* KEEP = "TRUE" *) wire n517;
    (* KEEP = "TRUE" *) wire n518;
    (* KEEP = "TRUE" *) wire n519;
    (* KEEP = "TRUE" *) wire n520;
    (* KEEP = "TRUE" *) wire n521;
    (* KEEP = "TRUE" *) wire n522;
    (* KEEP = "TRUE" *) wire n523;
    (* KEEP = "TRUE" *) wire n524;
    (* KEEP = "TRUE" *) wire n525;
    (* KEEP = "TRUE" *) wire n526;
    (* KEEP = "TRUE" *) wire n527;
    (* KEEP = "TRUE" *) wire n528;
    (* KEEP = "TRUE" *) wire n529;
    (* KEEP = "TRUE" *) wire n530;
    (* KEEP = "TRUE" *) wire n531;
    (* KEEP = "TRUE" *) wire n532;
    (* KEEP = "TRUE" *) wire n533;
    (* KEEP = "TRUE" *) wire n534;
    (* KEEP = "TRUE" *) wire n535;
    (* KEEP = "TRUE" *) wire n536;
    (* KEEP = "TRUE" *) wire n537;
    (* KEEP = "TRUE" *) wire n538;
    (* KEEP = "TRUE" *) wire n539;
    (* KEEP = "TRUE" *) wire n540;
    (* KEEP = "TRUE" *) wire n541;
    (* KEEP = "TRUE" *) wire n542;
    (* KEEP = "TRUE" *) wire n543;
    (* KEEP = "TRUE" *) wire n544;
    (* KEEP = "TRUE" *) wire n545;
    (* KEEP = "TRUE" *) wire n546;
    (* KEEP = "TRUE" *) wire n547;
    (* KEEP = "TRUE" *) wire n548;
    (* KEEP = "TRUE" *) wire n549;
    (* KEEP = "TRUE" *) wire n550;
    (* KEEP = "TRUE" *) wire n551;
    (* KEEP = "TRUE" *) wire n552;
    (* KEEP = "TRUE" *) wire n553;
    (* KEEP = "TRUE" *) wire n554;
    (* KEEP = "TRUE" *) wire n555;
    (* KEEP = "TRUE" *) wire n556;
    (* KEEP = "TRUE" *) wire n557;
    (* KEEP = "TRUE" *) wire n558;
    (* KEEP = "TRUE" *) wire n559;
    (* KEEP = "TRUE" *) wire n560;
    (* KEEP = "TRUE" *) wire n561;
    (* KEEP = "TRUE" *) wire n562;
    (* KEEP = "TRUE" *) wire n563;
    (* KEEP = "TRUE" *) wire n564;
    (* KEEP = "TRUE" *) wire n565;
    (* KEEP = "TRUE" *) wire n566;
    (* KEEP = "TRUE" *) wire n567;
    (* KEEP = "TRUE" *) wire n568;
    (* KEEP = "TRUE" *) wire n569;
    (* KEEP = "TRUE" *) wire n570;
    (* KEEP = "TRUE" *) wire n571;
    (* KEEP = "TRUE" *) wire n572;
    (* KEEP = "TRUE" *) wire n573;
    (* KEEP = "TRUE" *) wire n574;
    (* KEEP = "TRUE" *) wire n575;
    (* KEEP = "TRUE" *) wire n576;
    (* KEEP = "TRUE" *) wire n577;
    (* KEEP = "TRUE" *) wire n578;
    (* KEEP = "TRUE" *) wire n579;
    (* KEEP = "TRUE" *) wire n580;
    (* KEEP = "TRUE" *) wire n581;
    (* KEEP = "TRUE" *) wire n582;
    (* KEEP = "TRUE" *) wire n583;
    (* KEEP = "TRUE" *) wire n584;
    (* KEEP = "TRUE" *) wire n585;
    (* KEEP = "TRUE" *) wire n586;
    (* KEEP = "TRUE" *) wire n587;
    (* KEEP = "TRUE" *) wire n588;
    (* KEEP = "TRUE" *) wire n589;
    (* KEEP = "TRUE" *) wire n590;
    (* KEEP = "TRUE" *) wire n591;
    (* KEEP = "TRUE" *) wire n592;
    (* KEEP = "TRUE" *) wire n593;
    (* KEEP = "TRUE" *) wire n594;
    (* KEEP = "TRUE" *) wire n595;
    (* KEEP = "TRUE" *) wire n596;
    (* KEEP = "TRUE" *) wire n597;
    (* KEEP = "TRUE" *) wire n598;
    (* KEEP = "TRUE" *) wire n599;
    (* KEEP = "TRUE" *) wire n600;
    (* KEEP = "TRUE" *) wire n601;
    (* KEEP = "TRUE" *) wire n602;
    (* KEEP = "TRUE" *) wire n603;
    (* KEEP = "TRUE" *) wire n604;
    (* KEEP = "TRUE" *) wire n605;
    (* KEEP = "TRUE" *) wire n606;
    (* KEEP = "TRUE" *) wire n607;
    (* KEEP = "TRUE" *) wire n608;
    (* KEEP = "TRUE" *) wire n609;
    (* KEEP = "TRUE" *) wire n610;
    (* KEEP = "TRUE" *) wire n611;
    (* KEEP = "TRUE" *) wire n612;
    (* KEEP = "TRUE" *) wire n613;
    (* KEEP = "TRUE" *) wire n614;
    (* KEEP = "TRUE" *) wire n615;
    (* KEEP = "TRUE" *) wire n616;
    (* KEEP = "TRUE" *) wire n617;
    (* KEEP = "TRUE" *) wire n618;
    (* KEEP = "TRUE" *) wire n619;
    (* KEEP = "TRUE" *) wire n620;
    (* KEEP = "TRUE" *) wire n621;
    (* KEEP = "TRUE" *) wire n622;
    (* KEEP = "TRUE" *) wire n623;
    (* KEEP = "TRUE" *) wire n624;
    (* KEEP = "TRUE" *) wire n625;
    (* KEEP = "TRUE" *) wire n626;
    (* KEEP = "TRUE" *) wire n627;
    (* KEEP = "TRUE" *) wire n628;
    (* KEEP = "TRUE" *) wire n629;
    (* KEEP = "TRUE" *) wire n630;
    (* KEEP = "TRUE" *) wire n631;
    (* KEEP = "TRUE" *) wire n632;
    (* KEEP = "TRUE" *) wire n633;
    (* KEEP = "TRUE" *) wire n634;
    (* KEEP = "TRUE" *) wire n635;
    (* KEEP = "TRUE" *) wire n636;
    (* KEEP = "TRUE" *) wire n637;
    (* KEEP = "TRUE" *) wire n638;
    (* KEEP = "TRUE" *) wire n639;
    (* KEEP = "TRUE" *) wire n640;
    (* KEEP = "TRUE" *) wire n641;
    (* KEEP = "TRUE" *) wire n642;
    (* KEEP = "TRUE" *) wire n643;
    (* KEEP = "TRUE" *) wire n644;
    (* KEEP = "TRUE" *) wire n645;
    (* KEEP = "TRUE" *) wire n646;
    (* KEEP = "TRUE" *) wire n647;
    (* KEEP = "TRUE" *) wire n648;
    (* KEEP = "TRUE" *) wire n649;
    (* KEEP = "TRUE" *) wire n650;
    (* KEEP = "TRUE" *) wire n651;
    (* KEEP = "TRUE" *) wire n652;

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5B0F4AD01917683C)) n0_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n0)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5A5A52F47776E968)) n1_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n1)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h02AAAAA2AE7777E8)) n2_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n2)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5400000471888815)) n3_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n3)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n4_lut (
        .I0(n0), .I1(n1), .I2(n2), .I3(n3), .I4(x[3]), .I5(x[9]), .O(n4)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h02020055869E7199)) n5_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n5)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBFFDFDBF9E8699E6)) n6_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n6)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBDF5F5FD1E87871E)) n7_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n7)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2FBDF5F578968796)) n8_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n8)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n9_lut (
        .I0(n5), .I1(n6), .I2(n7), .I3(n8), .I4(x[5]), .I5(x[9]), .O(n9)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h855E87E97887E761)) n10_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n10)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5FF8A15E6186799E)) n11_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n11)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBDD0BDD4F5AFFF0A)) n12_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n12)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD00B4A2F40D40A50)) n13_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n13)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n14_lut (
        .I0(n10), .I1(n11), .I2(n12), .I3(n13), .I4(x[6]), .I5(x[11]), .O(n14)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1FE817A11E617918)) n15_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n15)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE88107E879E79EE7)) n16_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n16)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD00B420B0A402A50)) n17_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n17)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4BBDBDF4BDAFD4BF)) n18_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n18)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n19_lut (
        .I0(n15), .I1(n16), .I2(n17), .I3(n18), .I4(x[6]), .I5(x[11]), .O(n19)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n20_lut (
        .I0(n4), .I1(n9), .I2(n14), .I3(n19), .I4(x[4]), .I5(x[8]), .O(n20)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE6E6E6869879E699)) n21_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n21)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE178785A5A7879E1)) n22_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n22)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2A54AB54AAD500BF)) n23_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n23)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2FBFBDFDF5F5FDBD)) n24_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n24)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n25_lut (
        .I0(n21), .I1(n22), .I2(n23), .I3(n24), .I4(x[9]), .I5(x[11]), .O(n25)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFDFFAA1939E663)) n26_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n26)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4002005039196198)) n27_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n27)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h50420A42E17A5861)) n28_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n28)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD4420A0285785A78)) n29_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n29)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n30_lut (
        .I0(n26), .I1(n27), .I2(n28), .I3(n29), .I4(x[5]), .I5(x[9]), .O(n30)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5EE15A87E5189E86)) n31_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n31)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE8851EA18618E779)) n32_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n32)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h520B420B025040F5)) n33_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n33)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0BB5BDD4AF2BFDAB)) n34_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n34)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n35_lut (
        .I0(n31), .I1(n32), .I2(n33), .I3(n34), .I4(x[6]), .I5(x[11]), .O(n35)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE887781E7986E761)) n36_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n36)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h055E7A87A79E799E)) n37_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n37)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2BB52FBDF5BFF5AB)) n38_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n38)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBDD2D00B40D42A40)) n39_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n39)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n40_lut (
        .I0(n36), .I1(n37), .I2(n38), .I3(n39), .I4(x[6]), .I5(x[11]), .O(n40)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n41_lut (
        .I0(n25), .I1(n30), .I2(n35), .I3(n40), .I4(x[4]), .I5(x[8]), .O(n41)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F0F18F300888813)) n42_lut (
        .I0(x[2]), .I1(x[3]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n42)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC1E30F30CEFFEEC8)) n43_lut (
        .I0(x[2]), .I1(x[3]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n43)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h83C38F18EF7777FE)) n44_lut (
        .I0(x[2]), .I1(x[3]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n44)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0F0F18F73100137)) n45_lut (
        .I0(x[2]), .I1(x[3]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n45)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n46_lut (
        .I0(n42), .I1(n43), .I2(n44), .I3(n45), .I4(x[0]), .I5(x[4]), .O(n46)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFEAAA000555FF)) n47_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n47)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000155555)) n48_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n48)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00AAABFFFF555554)) n49_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n49)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n50_lut (
        .I0(n47), .I1(n48), .I2(1'b0), .I3(n49), .I4(x[7]), .I5(x[8]), .O(n50)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB42DD4BDD0BDF42D)) n51_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[7]), .O(n51)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h42D00B422F422B42)) n52_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[7]), .O(n52)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC2D2BC2D42D22D0B)) n53_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[7]), .O(n53)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4B4BD0B42F4BF4BD)) n54_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[7]), .O(n54)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n55_lut (
        .I0(n51), .I1(n52), .I2(n53), .I3(n54), .I4(x[5]), .I5(x[8]), .O(n55)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0AFF54000000015F)) n56_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n56)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h502BFFD555555FFE)) n57_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n57)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF500AAFFFFFFFFA8)) n58_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n58)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hAFD5002AAAAAA800)) n59_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n59)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n60_lut (
        .I0(n56), .I1(n57), .I2(n58), .I3(n59), .I4(x[2]), .I5(x[3]), .O(n60)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n61_lut (
        .I0(n46), .I1(n50), .I2(n55), .I3(n60), .I4(x[9]), .I5(x[11]), .O(n61)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF870F58AF75557FE)) n62_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n62)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5A5A70AF51000157)) n63_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n63)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5E1A58F518AAAA81)) n64_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n64)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1F0F1A718AEFFFEA)) n65_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n65)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n66_lut (
        .I0(n62), .I1(n63), .I2(n64), .I3(n65), .I4(x[3]), .I5(x[4]), .O(n66)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h80001555FFFEAA00)) n67_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n67)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF555500002AAAAA)) n68_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n68)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n69_lut (
        .I0(n67), .I1(~(n48)), .I2(1'b1), .I3(n68), .I4(x[7]), .I5(x[8]), .O(n69)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBB20B2044DB24DB0)) n70_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n70)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h44DD4DDBB20DF24D)) n71_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n71)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCDDF4CDFDB204DB2)) n72_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n72)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB220FB20204DFA05)) n73_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n73)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n74_lut (
        .I0(n70), .I1(n71), .I2(n72), .I3(n73), .I4(x[3]), .I5(x[6]), .O(n74)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4022223322220044)) n75_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n75)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBBFDDDDCCDDDDFBB)) n76_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n76)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3BBDDCC433BBB333)) n77_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n77)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hDC40223BCC4444CC)) n78_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n78)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n79_lut (
        .I0(n75), .I1(n76), .I2(n77), .I3(n78), .I4(x[3]), .I5(x[7]), .O(n79)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n80_lut (
        .I0(n66), .I1(n69), .I2(n74), .I3(n79), .I4(x[9]), .I5(x[11]), .O(n80)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n81_lut (
        .I0(n20), .I1(n41), .I2(n61), .I3(n80), .I4(x[1]), .I5(x[10]), .O(n81)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8C7388FFC1C31778)) n82_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n82)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEF8C10F7837C17C1)) n83_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n83)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF7F7F7EC7CFCE8)) n84_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n84)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF7108CEF37E817C1)) n85_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n85)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n86_lut (
        .I0(n82), .I1(n83), .I2(n84), .I3(n85), .I4(x[8]), .I5(x[9]), .O(n86)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h78EE0F7EFE371771)) n87_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n87)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0CC0EFE3701C11E)) n88_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n88)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE0EEC3001073CC7E)) n89_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n89)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h838C83008C187783)) n90_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n90)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n91_lut (
        .I0(n87), .I1(n88), .I2(n89), .I3(n90), .I4(x[3]), .I5(x[6]), .O(n91)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC8FC7CE83E3E7CC3)) n92_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[9]), .O(n92)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEC817E83C137C17C)) n93_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[9]), .O(n93)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1008080811EF10CE)) n94_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[9]), .O(n94)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h108EF7310031F7CC)) n95_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[9]), .O(n95)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n96_lut (
        .I0(n92), .I1(n93), .I2(n94), .I3(n95), .I4(x[8]), .I5(x[11]), .O(n96)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4FDDF020887781C3)) n97_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n97)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F00D2FBFF00EC68)) n98_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n98)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF2FDDBFDF3F3E789)) n99_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n99)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hDB400F00101831EE)) n100_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n100)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n101_lut (
        .I0(n97), .I1(n98), .I2(n99), .I3(n100), .I4(x[1]), .I5(x[6]), .O(n101)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n102_lut (
        .I0(n86), .I1(n91), .I2(n96), .I3(n101), .I4(x[4]), .I5(x[5]), .O(n102)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7E817C133C1683C3)) n103_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n103)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC813C03717C17C17)) n104_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n104)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7100731000881110)) n105_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n105)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h08CFFF31EF731008)) n106_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n106)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n107_lut (
        .I0(n103), .I1(n104), .I2(n105), .I3(n106), .I4(x[8]), .I5(x[11]), .O(n107)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF773733317C13E17)) n108_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[8]), .I5(x[11]), .O(n108)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h08CE331083E8C1E8)) n109_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[8]), .I5(x[11]), .O(n109)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h108CCEFF817E7E83)) n110_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[8]), .I5(x[11]), .O(n110)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCF738CFF037E7E81)) n111_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[8]), .I5(x[11]), .O(n111)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n112_lut (
        .I0(n108), .I1(n109), .I2(n110), .I3(n111), .I4(x[7]), .I5(x[9]), .O(n112)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h31EF77F73E7C177C)) n113_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n113)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF78CFFFFC1C13EE8)) n114_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n114)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h08F71008C8EC8381)) n115_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n115)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF3CE73317F37FC7E)) n116_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n116)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n117_lut (
        .I0(n113), .I1(n114), .I2(n115), .I3(n116), .I4(x[4]), .I5(x[9]), .O(n117)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h10F700EEC08117C1)) n118_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n118)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF3CE31CC7E7E7C83)) n119_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n119)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCFEFEFEE131317E8)) n120_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n120)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h10088C8CC8E8E8C3)) n121_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[8]), .I4(x[9]), .I5(x[11]), .O(n121)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n122_lut (
        .I0(n118), .I1(n119), .I2(n120), .I3(n121), .I4(x[4]), .I5(x[7]), .O(n122)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n123_lut (
        .I0(n107), .I1(n112), .I2(n117), .I3(n122), .I4(x[5]), .I5(x[6]), .O(n123)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1137EC80137EC801)) n124_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n124)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h33337777FFFEEECC)) n125_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n125)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF308EF710CF7308E)) n126_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n126)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h308F708E710EF30C)) n127_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n127)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n128_lut (
        .I0(n124), .I1(n125), .I2(n126), .I3(n127), .I4(x[9]), .I5(x[11]), .O(n128)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h377FEC801337EEC8)) n129_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n129)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000111111)) n130_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n130)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF710CF710CF7108E)) n131_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n131)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h30CF30CF30CF30CF)) n132_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n132)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n133_lut (
        .I0(n129), .I1(n130), .I2(n131), .I3(n132), .I4(x[9]), .I5(x[11]), .O(n133)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h88011337FEEC8801)) n134_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n134)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0CF308EF308E710C)) n135_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n135)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF10EF18F708F70CF)) n136_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n136)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n137_lut (
        .I0(n134), .I1(1'b0), .I2(n135), .I3(n136), .I4(x[9]), .I5(x[11]), .O(n137)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7733111080137FEC)) n138_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n138)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF773311880137FE)) n139_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n139)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h30180C0C08103071)) n140_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n140)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8FEFF7F3F3F7EF8F)) n141_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n141)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n142_lut (
        .I0(n138), .I1(n139), .I2(n140), .I3(n141), .I4(x[4]), .I5(x[11]), .O(n142)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n143_lut (
        .I0(n128), .I1(n133), .I2(n137), .I3(n142), .I4(x[7]), .I5(x[8]), .O(n143)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCC880133C837807E)) n144_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n144)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFEEE8037C837)) n145_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n145)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF7FC813FE)) n146_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n146)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h88CCEEEE7FEE8813)) n147_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n147)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n148_lut (
        .I0(n144), .I1(n145), .I2(n146), .I3(n147), .I4(x[7]), .I5(x[8]), .O(n148)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCCC80011FE01EC13)) n149_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n149)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFEEEC13FE01)) n150_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n150)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF37EE8037)) n151_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n151)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0088CCEE37FECC01)) n152_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n152)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n153_lut (
        .I0(n149), .I1(n150), .I2(n151), .I3(n152), .I4(x[7]), .I5(x[8]), .O(n153)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFEC0037FC03FC03)) n154_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n154)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEC8013FFC01FE81F)) n155_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n155)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEFF7331111111337)) n156_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n156)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0CEEFFFFF77FFFFF)) n157_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n157)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n158_lut (
        .I0(n154), .I1(n155), .I2(n156), .I3(n157), .I4(x[3]), .I5(x[9]), .O(n158)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00037FEC017E807E)) n159_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n159)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h137FFE8017FC03F8)) n160_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n160)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h10008CCEEEEEECC8)) n161_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n161)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF731000008800000)) n162_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n162)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n163_lut (
        .I0(n159), .I1(n160), .I2(n161), .I3(n162), .I4(x[3]), .I5(x[9]), .O(n163)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n164_lut (
        .I0(n148), .I1(n153), .I2(n158), .I3(n163), .I4(x[4]), .I5(x[11]), .O(n164)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n165_lut (
        .I0(n102), .I1(n123), .I2(n143), .I3(n164), .I4(x[2]), .I5(x[10]), .O(n165)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFE3FFE077E3EC0)) n166_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[8]), .I5(x[10]), .O(n166)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F3F030F7EE0FC83)) n167_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[8]), .I5(x[10]), .O(n167)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0307E080E007F007)) n168_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[8]), .I5(x[10]), .O(n168)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8001FEF8077EC11F)) n169_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[8]), .I5(x[10]), .O(n169)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n170_lut (
        .I0(n166), .I1(n167), .I2(n168), .I3(n169), .I4(x[5]), .I5(x[6]), .O(n170)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h03071F7F1FF0077C)) n171_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n171)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8F0C080C00FF881)) n172_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n172)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8F0E0C0C0077EE0)) n173_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n173)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFFFEFCF0811FFC)) n174_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n174)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n175_lut (
        .I0(n171), .I1(n172), .I2(n173), .I3(n174), .I4(x[6]), .I5(x[8]), .O(n175)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFEFF1FFCFF7FFFF)) n176_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n176)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0F700F3FF00F710)) n177_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n177)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0C00CF0808FFEFFF)) n178_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n178)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8F0CFF8FEF73FF33)) n179_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n179)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n180_lut (
        .I0(n176), .I1(n177), .I2(n178), .I3(n179), .I4(x[2]), .I5(x[5]), .O(n180)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7F0700C0C0F0F8FC)) n181_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n181)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0700E0FE03010080)) n182_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n182)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0FF3F01070100C0)) n183_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n183)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFCFF0700FEFF7F1F)) n184_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n184)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n185_lut (
        .I0(n181), .I1(n182), .I2(n183), .I3(n184), .I4(x[6]), .I5(x[8]), .O(n185)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n186_lut (
        .I0(n170), .I1(n175), .I2(n180), .I3(n185), .I4(x[7]), .I5(x[11]), .O(n186)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0FF8037EC01FF007)) n187_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n187)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h01030F3FFEF8E080)) n188_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n188)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0301000080C0E0E0)) n189_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n189)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F00C0F8FF1F0300)) n190_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n190)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n191_lut (
        .I0(n187), .I1(n188), .I2(n189), .I3(n190), .I4(x[10]), .I5(x[11]), .O(n191)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFEFCF0C0F8033EE0)) n192_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n192)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h03071F3F0FFCC01F)) n193_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n193)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00E0FEFF3F1F0F07)) n194_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n194)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE0FE7F07FCFEFF7F)) n195_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n195)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n196_lut (
        .I0(n192), .I1(n193), .I2(n194), .I3(n195), .I4(x[6]), .I5(x[11]), .O(n196)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0301E0F0077E7EE0)) n197_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n197)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3F0F00807EE0E007)) n198_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n198)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00C00700FEFCC000)) n199_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n199)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF1FFCFF3F7FF0E0)) n200_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n200)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n201_lut (
        .I0(n197), .I1(n198), .I2(n199), .I3(n200), .I4(x[5]), .I5(x[10]), .O(n201)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0FCFF7F0FFCE007)) n202_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[11]), .O(n202)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h030000C0031FF8C0)) n203_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[11]), .O(n203)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7F0300F803070F1F)) n204_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[11]), .O(n204)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1F00C0FEC0800001)) n205_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[11]), .O(n205)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n206_lut (
        .I0(n202), .I1(n203), .I2(n204), .I3(n205), .I4(x[6]), .I5(x[10]), .O(n206)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n207_lut (
        .I0(n191), .I1(n196), .I2(n201), .I3(n206), .I4(x[7]), .I5(x[8]), .O(n207)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1700F8FE7F3F3F7F)) n208_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n208)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FC7F0703010103)) n209_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n209)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h80FE3F0380C0C0C0)) n210_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n210)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC3F00E0FCFEFEFC)) n211_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n211)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n212_lut (
        .I0(n208), .I1(n209), .I2(n210), .I3(n211), .I4(x[2]), .I5(x[5]), .O(n212)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h030307070F1F1F3F)) n213_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n213)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000010101)) n214_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n214)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F07070303010100)) n215_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n215)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n216_lut (
        .I0(n213), .I1(n214), .I2(1'b0), .I3(n215), .I4(x[7]), .I5(x[8]), .O(n216)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0100E0F80100C0F8)) n217_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n217)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFCFF3F0FFE7F1F07)) n218_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n218)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF3F07000F0100E0)) n219_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n219)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0700C0F8C0F8FF7F)) n220_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n220)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n221_lut (
        .I0(n217), .I1(n218), .I2(n219), .I3(n220), .I4(x[6]), .I5(x[8]), .O(n221)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF030100000000030)) n222_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n222)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00080C0E0E0E0C08)) n223_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n223)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F8FEFFFFFFFFFEF)) n224_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n224)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEFFFF3F1F1F1F1F3)) n225_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n225)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n226_lut (
        .I0(n222), .I1(n223), .I2(n224), .I3(n225), .I4(x[2]), .I5(x[5]), .O(n226)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n227_lut (
        .I0(n212), .I1(n216), .I2(n221), .I3(n226), .I4(x[10]), .I5(x[11]), .O(n227)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC3F0180E0F8F0E0)) n228_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n228)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7F01C0FCFF7F7F7E)) n229_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n229)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3F00F8FF3F1F071F)) n230_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n230)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h01F87F0701808080)) n231_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n231)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n232_lut (
        .I0(n228), .I1(n229), .I2(n230), .I3(n231), .I4(x[2]), .I5(x[5]), .O(n232)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h002AFFFFFFEA0000)) n233_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n233)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2BFFFFFFFFFFFA00)) n234_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n234)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFFF8)) n235_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n235)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n236_lut (
        .I0(n233), .I1(n234), .I2(n235), .I3(1'b1), .I4(x[1]), .I5(x[2]), .O(n236)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFCFF7F0FFCFF7F1F)) n237_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n237)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h070180E00300C0F0)) n238_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n238)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0180F0FEE0FCFF3F)) n239_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n239)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE0FEFF0FFF1F0300)) n240_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[7]), .O(n240)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n241_lut (
        .I0(n237), .I1(n238), .I2(n239), .I3(n240), .I4(x[6]), .I5(x[8]), .O(n241)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFEFFFFFF7FFFFFFF)) n242_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n242)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h80E0F0F8FCFCF8F0)) n243_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n243)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0300000000800000)) n244_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n244)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF3F0F0703030307)) n245_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n245)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n246_lut (
        .I0(n242), .I1(n243), .I2(n244), .I3(n245), .I4(x[4]), .I5(x[5]), .O(n246)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n247_lut (
        .I0(n232), .I1(n236), .I2(n241), .I3(n246), .I4(x[10]), .I5(x[11]), .O(n247)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n248_lut (
        .I0(n186), .I1(n207), .I2(n227), .I3(n247), .I4(x[3]), .I5(x[9]), .O(n248)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00C03F0FF000FC00)) n249_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[10]), .I5(x[11]), .O(n249)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF01FF7FFFFFE007)) n250_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[10]), .I5(x[11]), .O(n250)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF7FC0F8C000FF80)) n251_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[10]), .I5(x[11]), .O(n251)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00F00000FEF88007)) n252_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[10]), .I5(x[11]), .O(n252)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n253_lut (
        .I0(n249), .I1(n250), .I2(n251), .I3(n252), .I4(x[6]), .I5(x[8]), .O(n253)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h033FFFFFFF801FF8)) n254_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n254)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFFFFFFFF8007FF)) n255_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n255)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000E0FF01000000)) n256_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n256)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE0FFFF00F0FEFFFF)) n257_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n257)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n258_lut (
        .I0(n254), .I1(n255), .I2(n256), .I3(n257), .I4(x[8]), .I5(x[11]), .O(n258)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFEFFFFFF0FFE007F)) n259_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n259)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF1F0100FE0007FF)) n260_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n260)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000F8FF0000077F)) n261_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n261)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FFFF01FFFFFFFF)) n262_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n262)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n263_lut (
        .I0(n259), .I1(n260), .I2(n261), .I3(n262), .I4(x[8]), .I5(x[10]), .O(n263)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8C00000001FFC00)) n264_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n264)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0001071F1FFF0007)) n265_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n265)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00F8FFFFFF7F1F07)) n266_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n266)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF030000000080)) n267_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n267)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n268_lut (
        .I0(n264), .I1(n265), .I2(n266), .I3(n267), .I4(x[8]), .I5(x[11]), .O(n268)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n269_lut (
        .I0(n253), .I1(n258), .I2(n263), .I3(n268), .I4(x[3]), .I5(x[7]), .O(n269)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h037F003FFF07FF3F)) n270_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n270)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000F00007800300)) n271_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n271)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000F000307800100)) n272_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n272)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC000FE0080FFF0FF)) n273_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n273)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n274_lut (
        .I0(n270), .I1(n271), .I2(n272), .I3(n273), .I4(x[3]), .I5(x[5]), .O(n274)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFCE0FF001FF8)) n275_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n275)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h031FFFFF0FFF003F)) n276_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n276)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h80000000001FFF80)) n277_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n277)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFCF0FC000FFF)) n278_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n278)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n279_lut (
        .I0(n275), .I1(n276), .I2(n277), .I3(n278), .I4(x[3]), .I5(x[8]), .O(n279)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF03FFFFC0FFE0)) n280_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n280)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF000FFF0FC00FF00)) n281_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n281)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000F800007F000F)) n282_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n282)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00FF3FFF03FF)) n283_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n283)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n284_lut (
        .I0(n280), .I1(n281), .I2(n282), .I3(n283), .I4(x[6]), .I5(x[8]), .O(n284)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00030000C000F000)) n285_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n285)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC00FF80FFF8FFFF)) n286_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n286)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF87FFF007F0000)) n287_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n287)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1FFF00078000FFC0)) n288_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n288)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n289_lut (
        .I0(n285), .I1(n286), .I2(n287), .I3(n288), .I4(x[8]), .I5(x[10]), .O(n289)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n290_lut (
        .I0(n274), .I1(n279), .I2(n284), .I3(n289), .I4(x[7]), .I5(x[11]), .O(n290)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF037F001F003F)) n291_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n291)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h001F8000F000F000)) n292_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n292)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0007F000FFC0FFE0)) n293_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n293)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE000FFFE1FFF07FF)) n294_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n294)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n295_lut (
        .I0(n291), .I1(n292), .I2(n293), .I3(n294), .I4(x[3]), .I5(x[6]), .O(n295)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h73100000001137FF)) n296_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n296)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000000013)) n297_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n297)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n298_lut (
        .I0(n296), .I1(n297), .I2(1'b0), .I3(1'b0), .I4(x[2]), .I5(x[3]), .O(n298)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFE3FFFFFFF1FFF)) n299_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n299)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE000FF80FF80FFF8)) n300_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n300)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h003F00000000F000)) n301_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n301)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0FFF01FF000F)) n302_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n302)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n303_lut (
        .I0(n299), .I1(n300), .I2(n301), .I3(n302), .I4(x[6]), .I5(x[7]), .O(n303)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FF001F001F003F)) n304_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n304)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF7FFFFFFF)) n305_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n305)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC00FFC0FFE0FFE0)) n306_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n306)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n307_lut (
        .I0(1'b0), .I1(n304), .I2(n305), .I3(n306), .I4(x[5]), .I5(x[6]), .O(n307)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n308_lut (
        .I0(n295), .I1(n298), .I2(n303), .I3(n307), .I4(x[10]), .I5(x[11]), .O(n308)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h01FF7FFC01FF7FF8)) n309_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n309)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC000007FF008003)) n310_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n310)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFC0FC000FFFFFF0)) n311_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n311)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h03FF7FFE8003007F)) n312_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n312)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n313_lut (
        .I0(n309), .I1(n310), .I2(n311), .I3(n312), .I4(x[6]), .I5(x[8]), .O(n313)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h08CEFFFFFFFEC800)) n314_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n314)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFFFE)) n315_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n315)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n316_lut (
        .I0(n314), .I1(n315), .I2(1'b1), .I3(1'b1), .I4(x[2]), .I5(x[3]), .O(n316)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000F000000018000)) n317_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n317)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF03FF03FF001F)) n318_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n318)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFE00FFF8FFFE7FFF)) n319_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n319)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00070000F800FFC0)) n320_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[8]), .O(n320)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n321_lut (
        .I0(n317), .I1(n318), .I2(n319), .I3(n320), .I4(x[6]), .I5(x[7]), .O(n321)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFCFFFFFFFFFFFC)) n322_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n322)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC000F800FC00F800)) n323_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n323)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000F000100000000)) n324_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n324)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0FFF03FF03FF)) n325_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n325)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n326_lut (
        .I0(n322), .I1(n323), .I2(n324), .I3(n325), .I4(x[5]), .I5(x[6]), .O(n326)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n327_lut (
        .I0(n313), .I1(n316), .I2(n321), .I3(n326), .I4(x[10]), .I5(x[11]), .O(n327)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n328_lut (
        .I0(n269), .I1(n290), .I2(n308), .I3(n327), .I4(x[4]), .I5(x[9]), .O(n328)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF80FFF0FFF80000)) n329_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n329)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF03FFFFC0)) n330_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n330)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFEFFFF3FFFFFFF)) n331_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n331)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF03FF0000003F)) n332_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n332)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n333_lut (
        .I0(n329), .I1(n330), .I2(n331), .I3(n332), .I4(x[4]), .I5(x[10]), .O(n333)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8000F800E000007F)) n334_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n334)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFC000)) n335_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n335)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000007F)) n336_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n336)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8000FFFFE0000000)) n337_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n337)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n338_lut (
        .I0(n334), .I1(n335), .I2(n336), .I3(n337), .I4(x[4]), .I5(x[10]), .O(n338)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF000000007FFFF)) n339_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n339)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC000000F8000007)) n340_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n340)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000007FFF800000)) n341_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n341)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FFFFFFFFFC0000)) n342_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n342)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n343_lut (
        .I0(n339), .I1(n340), .I2(n341), .I3(n342), .I4(x[6]), .I5(x[10]), .O(n343)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h001F0000FFFFF800)) n344_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n344)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000001FFFFF)) n345_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n345)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFEFE00E000)) n346_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n346)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF8FFFFFFFFFFFF)) n347_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[11]), .O(n347)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n348_lut (
        .I0(n344), .I1(n345), .I2(n346), .I3(n347), .I4(x[4]), .I5(x[10]), .O(n348)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n349_lut (
        .I0(n333), .I1(n338), .I2(n343), .I3(n348), .I4(x[7]), .I5(x[8]), .O(n349)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC00000000001FFF)) n350_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n350)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFCFFFE0000)) n351_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n351)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFFFFFFFFFFF800)) n352_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n352)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000F0007FFFF)) n353_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n353)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n354_lut (
        .I0(n350), .I1(n351), .I2(n352), .I3(n353), .I4(x[4]), .I5(x[8]), .O(n354)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF000000F001FFFFF)) n355_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n355)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFE000F0000007)) n356_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n356)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h03FFFFFFFFFFFFF8)) n357_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n357)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000FF000007FF)) n358_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n358)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n359_lut (
        .I0(n355), .I1(n356), .I2(n357), .I3(n358), .I4(x[8]), .I5(x[10]), .O(n359)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000001FF0000003F)) n360_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n360)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3FFFFFFF007FFFFF)) n361_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n361)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000FF00000000)) n362_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n362)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFF0000)) n363_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n363)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n364_lut (
        .I0(n360), .I1(n361), .I2(n362), .I3(n363), .I4(x[8]), .I5(x[10]), .O(n364)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFF1FFF)) n365_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n365)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF007F00030000)) n366_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n366)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF03FFFF00FFFE)) n367_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n367)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1FFF0000FFFFFFFF)) n368_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n368)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n369_lut (
        .I0(n365), .I1(n366), .I2(n367), .I3(n368), .I4(x[4]), .I5(x[8]), .O(n369)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n370_lut (
        .I0(n354), .I1(n359), .I2(n364), .I3(n369), .I4(x[7]), .I5(x[11]), .O(n370)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000007F0000003F)) n371_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n371)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF800000FFFC8000)) n372_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n372)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF8E000FFFFFFE0)) n373_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n373)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFFFFFF00077FFF)) n374_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n374)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n375_lut (
        .I0(n371), .I1(n372), .I2(n373), .I3(n374), .I4(x[4]), .I5(x[7]), .O(n375)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFCFFFFFFFFFEF8C0)) n376_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n376)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n377_lut (
        .I0(n376), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[3]), .I5(x[4]), .O(n377)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h001FFFFF00001FFF)) n378_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n378)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFF07FFFFFFF)) n379_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n379)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC000000FFFFC000)) n380_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n380)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000FFF00000000)) n381_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n381)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n382_lut (
        .I0(n378), .I1(n379), .I2(n380), .I3(n381), .I4(x[7]), .I5(x[8]), .O(n382)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0001FFFF0000FFFF)) n383_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n383)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF00000FFFF8000)) n384_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n384)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n385_lut (
        .I0(1'b0), .I1(n383), .I2(1'b1), .I3(n384), .I4(x[6]), .I5(x[7]), .O(n385)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n386_lut (
        .I0(n375), .I1(n377), .I2(n382), .I3(n385), .I4(x[10]), .I5(x[11]), .O(n386)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFC07FFFFFF)) n387_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n387)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00030FFF000001FF)) n388_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n388)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000FFE0000000)) n389_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n389)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC000000FFFFFE00)) n390_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[8]), .O(n390)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n391_lut (
        .I0(n387), .I1(n388), .I2(n389), .I3(n390), .I4(x[4]), .I5(x[7]), .O(n391)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h070100000001031F)) n392_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n392)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n393_lut (
        .I0(n392), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[3]), .I5(x[4]), .O(n393)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC000000FFFE0000)) n394_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n394)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000001FF00000000)) n395_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n395)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF000FFFFF)) n396_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n396)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF80000FFFFFFC0)) n397_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n397)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n398_lut (
        .I0(n394), .I1(n395), .I2(n396), .I3(n397), .I4(x[7]), .I5(x[8]), .O(n398)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFE0FFFFFFC0)) n399_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n399)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0000000FC000000)) n400_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n400)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000FF0000001F)) n401_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n401)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF03FFFFFF)) n402_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n402)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n403_lut (
        .I0(n399), .I1(n400), .I2(n401), .I3(n402), .I4(x[6]), .I5(x[7]), .O(n403)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n404_lut (
        .I0(n391), .I1(n393), .I2(n398), .I3(n403), .I4(x[10]), .I5(x[11]), .O(n404)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n405_lut (
        .I0(n349), .I1(n370), .I2(n386), .I3(n404), .I4(x[5]), .I5(x[9]), .O(n405)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0007FFFF00000000)) n406_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n406)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFFE000)) n407_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n407)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFFFF80)) n408_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n408)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFF8001FFFFF)) n409_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n409)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n410_lut (
        .I0(n406), .I1(n407), .I2(n408), .I3(n409), .I4(x[5]), .I5(x[7]), .O(n410)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFF80FFC00000)) n411_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n411)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000007FF000FFFFF)) n412_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n412)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n413_lut (
        .I0(n411), .I1(1'b1), .I2(1'b1), .I3(n412), .I4(x[5]), .I5(x[8]), .O(n413)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00001FFF0000003F)) n414_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n414)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF007FFFFF)) n415_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n415)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n416_lut (
        .I0(1'b1), .I1(n414), .I2(1'b1), .I3(n415), .I4(x[5]), .I5(x[8]), .O(n416)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF03FFFFFF)) n417_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n417)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h007FFFFF00000000)) n418_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n418)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFFFF80)) n419_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n419)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFC00FFFFFFFF)) n420_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n420)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n421_lut (
        .I0(n417), .I1(n418), .I2(n419), .I3(n420), .I4(x[5]), .I5(x[8]), .O(n421)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n422_lut (
        .I0(n410), .I1(n413), .I2(n416), .I3(n421), .I4(x[10]), .I5(x[11]), .O(n422)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFF803FFFFFF)) n423_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n423)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h001FFFFF00000000)) n424_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n424)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFFFFF0)) n425_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n425)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n426_lut (
        .I0(n423), .I1(n406), .I2(n424), .I3(n425), .I4(x[5]), .I5(x[7]), .O(n426)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000003FFF)) n427_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n427)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC00000000000000)) n428_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n428)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFF00FFFF8000)) n429_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n429)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n430_lut (
        .I0(n427), .I1(n428), .I2(1'b0), .I3(n429), .I4(x[5]), .I5(x[8]), .O(n430)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFC0000FFFFFE00)) n431_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n431)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000001F00000000)) n432_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n432)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000C0000000)) n433_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n433)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n434_lut (
        .I0(1'b0), .I1(n431), .I2(n432), .I3(n433), .I4(x[5]), .I5(x[8]), .O(n434)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFF0000000000)) n435_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n435)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000FFFFFF)) n436_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n436)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1FFFFFFFFFFFFFFF)) n437_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n437)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n438_lut (
        .I0(n435), .I1(1'b0), .I2(n436), .I3(n437), .I4(x[7]), .I5(x[8]), .O(n438)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n439_lut (
        .I0(n426), .I1(n430), .I2(n434), .I3(n438), .I4(x[10]), .I5(x[11]), .O(n439)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFFFFFFFFFFFFC0)) n440_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n440)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000007F)) n441_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n441)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n442_lut (
        .I0(n440), .I1(n441), .I2(1'b1), .I3(1'b1), .I4(x[8]), .I5(x[10]), .O(n442)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000001F01FFFFFF)) n443_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n443)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000100000000)) n444_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n444)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000F0000000)) n445_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n445)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000001FFFFFF00)) n446_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n446)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n447_lut (
        .I0(n443), .I1(n444), .I2(n445), .I3(n446), .I4(x[7]), .I5(x[8]), .O(n447)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFFE000)) n448_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n448)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF80000000)) n449_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n449)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF00000000)) n450_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[10]), .O(n450)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n451_lut (
        .I0(n448), .I1(n449), .I2(n450), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n451)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFF00000)) n452_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n452)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFF00FFFFFFFF)) n453_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n453)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n454_lut (
        .I0(1'b1), .I1(n452), .I2(n432), .I3(n453), .I4(x[8]), .I5(x[10]), .O(n454)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n455_lut (
        .I0(n442), .I1(n447), .I2(n451), .I3(n454), .I4(x[5]), .I5(x[11]), .O(n455)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF8000000000000)) n456_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n456)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFFFFFFFFFFFFFF)) n457_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n457)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF001FFFFF)) n458_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n458)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFF000FFFFFFFF)) n459_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n459)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n460_lut (
        .I0(n456), .I1(n457), .I2(n458), .I3(n459), .I4(x[8]), .I5(x[11]), .O(n460)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFF800)) n461_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n461)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000003FFFF)) n462_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n462)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000001FF00000000)) n463_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n463)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n464_lut (
        .I0(n461), .I1(n462), .I2(n463), .I3(1'b1), .I4(x[8]), .I5(x[11]), .O(n464)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFF0000)) n465_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n465)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF0001FFFF)) n466_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[7]), .O(n466)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n467_lut (
        .I0(1'b0), .I1(1'b0), .I2(n465), .I3(n466), .I4(x[8]), .I5(x[11]), .O(n467)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF8FFFFFFFFFFFC)) n468_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n468)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00000000FFFF)) n469_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n469)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0000FC00FFFF)) n470_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n470)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n471_lut (
        .I0(n468), .I1(1'b1), .I2(n469), .I3(n470), .I4(x[3]), .I5(x[11]), .O(n471)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n472_lut (
        .I0(n460), .I1(n464), .I2(n467), .I3(n471), .I4(x[5]), .I5(x[10]), .O(n472)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n473_lut (
        .I0(n422), .I1(n439), .I2(n455), .I3(n472), .I4(x[6]), .I5(x[9]), .O(n473)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00001FFFFFF80000)) n474_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n474)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n475_lut (
        .I0(1'b0), .I1(1'b0), .I2(n474), .I3(n474), .I4(x[0]), .I5(x[11]), .O(n475)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFF80000)) n476_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n476)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF0000000000000)) n477_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n477)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF80000000000000)) n478_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n478)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n479_lut (
        .I0(n476), .I1(n477), .I2(n478), .I3(1'b1), .I4(x[10]), .I5(x[11]), .O(n479)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h01FFFFFFFFFFFFFF)) n480_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n480)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFE000000000)) n481_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n481)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n482_lut (
        .I0(n480), .I1(n481), .I2(1'b0), .I3(1'b1), .I4(x[10]), .I5(x[11]), .O(n482)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000007F)) n483_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n483)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FFFFFFFF)) n484_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n484)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n485_lut (
        .I0(n483), .I1(1'b0), .I2(1'b0), .I3(n484), .I4(x[5]), .I5(x[10]), .O(n485)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n486_lut (
        .I0(n475), .I1(n479), .I2(n482), .I3(n485), .I4(x[8]), .I5(x[9]), .O(n486)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFC000000)) n487_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n487)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF0007FFFF)) n488_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[11]), .O(n488)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n489_lut (
        .I0(n487), .I1(1'b1), .I2(1'b1), .I3(n488), .I4(x[5]), .I5(x[8]), .O(n489)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFC000000000000)) n490_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n490)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFE00000)) n491_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n491)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n492_lut (
        .I0(1'b0), .I1(n490), .I2(n491), .I3(1'b0), .I4(x[8]), .I5(x[11]), .O(n492)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFC000)) n493_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n493)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FFFFFF00000000)) n494_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n494)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n495_lut (
        .I0(n493), .I1(1'b1), .I2(n494), .I3(1'b0), .I4(x[5]), .I5(x[11]), .O(n495)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFE0000)) n496_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n496)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n497_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(n496), .I4(x[8]), .I5(x[11]), .O(n497)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n498_lut (
        .I0(n489), .I1(n492), .I2(n495), .I3(n497), .I4(x[9]), .I5(x[10]), .O(n498)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h001FFFFFFFFFFFFF)) n499_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n499)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF80000000)) n500_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n500)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n501_lut (
        .I0(n499), .I1(1'b0), .I2(n500), .I3(1'b1), .I4(x[8]), .I5(x[9]), .O(n501)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000007FFFFFFFFFF)) n502_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n502)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000100000001)) n503_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[8]), .O(n503)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n504_lut (
        .I0(1'b1), .I1(n502), .I2(1'b1), .I3(n503), .I4(x[5]), .I5(x[9]), .O(n504)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00001FFFFFFFFFFF)) n505_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n505)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n506_lut (
        .I0(n505), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[8]), .I5(x[9]), .O(n506)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n507_lut (
        .I0(n478), .I1(1'b0), .I2(~(n481)), .I3(1'b1), .I4(x[8]), .I5(x[9]), .O(n507)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n508_lut (
        .I0(n501), .I1(n504), .I2(n506), .I3(n507), .I4(x[10]), .I5(x[11]), .O(n508)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n509_lut (
        .I0(1'b0), .I1(n491), .I2(1'b1), .I3(~(n500)), .I4(x[8]), .I5(x[9]), .O(n509)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n510_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[8]), .I5(x[9]), .O(n510)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000001F)) n511_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n511)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000001FFFFFFFFFF)) n512_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n512)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n513_lut (
        .I0(1'b0), .I1(n511), .I2(n512), .I3(1'b1), .I4(x[8]), .I5(x[9]), .O(n513)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n514_lut (
        .I0(1'b1), .I1(~(n437)), .I2(1'b0), .I3(1'b1), .I4(x[8]), .I5(x[9]), .O(n514)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n515_lut (
        .I0(n509), .I1(n510), .I2(n513), .I3(n514), .I4(x[10]), .I5(x[11]), .O(n515)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n516_lut (
        .I0(n486), .I1(n498), .I2(n508), .I3(n515), .I4(x[6]), .I5(x[7]), .O(n516)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n517_lut (
        .I0(1'b0), .I1(1'b0), .I2(~(n480)), .I3(1'b1), .I4(x[6]), .I5(x[9]), .O(n517)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n518_lut (
        .I0(~(n499)), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[9]), .O(n518)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n519_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[9]), .O(n519)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n520_lut (
        .I0(n505), .I1(1'b0), .I2(1'b1), .I3(n512), .I4(x[6]), .I5(x[9]), .O(n520)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n521_lut (
        .I0(n517), .I1(n518), .I2(n519), .I3(n520), .I4(x[7]), .I5(x[11]), .O(n521)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0007FFFFFFFFFFFF)) n522_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n522)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000007F)) n523_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n523)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n524_lut (
        .I0(1'b1), .I1(n522), .I2(n523), .I3(1'b0), .I4(x[6]), .I5(x[9]), .O(n524)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n525_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(n500), .I4(x[6]), .I5(x[9]), .O(n525)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n526_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[9]), .O(n526)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n527_lut (
        .I0(1'b0), .I1(~(n511)), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[9]), .O(n527)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n528_lut (
        .I0(n524), .I1(n525), .I2(n526), .I3(n527), .I4(x[7]), .I5(x[11]), .O(n528)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000001FFFFFFFF)) n529_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n529)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n530_lut (
        .I0(1'b1), .I1(1'b0), .I2(n529), .I3(1'b0), .I4(x[6]), .I5(x[9]), .O(n530)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFC000000)) n531_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n531)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n532_lut (
        .I0(n531), .I1(1'b1), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[9]), .O(n532)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n533_lut (
        .I0(1'b1), .I1(1'b1), .I2(n481), .I3(1'b1), .I4(x[6]), .I5(x[9]), .O(n533)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n534_lut (
        .I0(n519), .I1(n530), .I2(n532), .I3(n533), .I4(x[7]), .I5(x[11]), .O(n534)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFEFFFFF800)) n535_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[9]), .O(n535)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n536_lut (
        .I0(1'b0), .I1(n535), .I2(1'b1), .I3(1'b1), .I4(x[5]), .I5(x[6]), .O(n536)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n537_lut (
        .I0(1'b1), .I1(n436), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[9]), .O(n537)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n538_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[9]), .O(n538)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n539_lut (
        .I0(n526), .I1(n536), .I2(n537), .I3(n538), .I4(x[7]), .I5(x[11]), .O(n539)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n540_lut (
        .I0(n521), .I1(n528), .I2(n534), .I3(n539), .I4(x[8]), .I5(x[10]), .O(n540)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n541_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[10]), .I5(x[11]), .O(n541)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n542_lut (
        .I0(1'b0), .I1(1'b0), .I2(~(n505)), .I3(1'b0), .I4(x[10]), .I5(x[11]), .O(n542)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n543_lut (
        .I0(1'b0), .I1(1'b1), .I2(1'b1), .I3(1'b0), .I4(x[10]), .I5(x[11]), .O(n543)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n544_lut (
        .I0(n541), .I1(n541), .I2(n542), .I3(n543), .I4(x[6]), .I5(x[7]), .O(n544)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n545_lut (
        .I0(~(n522)), .I1(1'b1), .I2(1'b1), .I3(~(n436)), .I4(x[10]), .I5(x[11]), .O(n545)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n546_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[10]), .I5(x[11]), .O(n546)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n547_lut (
        .I0(n543), .I1(n545), .I2(n546), .I3(n546), .I4(x[6]), .I5(x[7]), .O(n547)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n548_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[7]), .O(n548)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n549_lut (
        .I0(1'b1), .I1(1'b1), .I2(n529), .I3(1'b0), .I4(x[6]), .I5(x[7]), .O(n549)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n550_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(n512), .I4(x[6]), .I5(x[7]), .O(n550)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n551_lut (
        .I0(n548), .I1(n549), .I2(n550), .I3(n548), .I4(x[10]), .I5(x[11]), .O(n551)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n552_lut (
        .I0(n523), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[7]), .O(n552)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n553_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[7]), .O(n553)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n554_lut (
        .I0(n552), .I1(n553), .I2(n553), .I3(n548), .I4(x[10]), .I5(x[11]), .O(n554)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n555_lut (
        .I0(n544), .I1(n547), .I2(n551), .I3(n554), .I4(x[8]), .I5(x[9]), .O(n555)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n556_lut (
        .I0(n553), .I1(n553), .I2(n553), .I3(n553), .I4(x[8]), .I5(x[11]), .O(n556)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n557_lut (
        .I0(~(n523)), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[7]), .O(n557)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n558_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(~(n512)), .I4(x[6]), .I5(x[7]), .O(n558)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n559_lut (
        .I0(n553), .I1(n557), .I2(n558), .I3(n548), .I4(x[8]), .I5(x[11]), .O(n559)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n560_lut (
        .I0(n548), .I1(n548), .I2(n548), .I3(n548), .I4(x[8]), .I5(x[11]), .O(n560)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n561_lut (
        .I0(n549), .I1(n553), .I2(n548), .I3(n548), .I4(x[8]), .I5(x[11]), .O(n561)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n562_lut (
        .I0(n556), .I1(n559), .I2(n560), .I3(n561), .I4(x[9]), .I5(x[10]), .O(n562)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n563_lut (
        .I0(n553), .I1(n553), .I2(n553), .I3(n553), .I4(x[8]), .I5(x[9]), .O(n563)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n564_lut (
        .I0(1'b0), .I1(1'b0), .I2(~(n529)), .I3(1'b1), .I4(x[6]), .I5(x[7]), .O(n564)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n565_lut (
        .I0(n553), .I1(n553), .I2(n564), .I3(n548), .I4(x[8]), .I5(x[9]), .O(n565)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n566_lut (
        .I0(n548), .I1(n548), .I2(n548), .I3(n548), .I4(x[8]), .I5(x[9]), .O(n566)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n567_lut (
        .I0(n563), .I1(n565), .I2(n566), .I3(n566), .I4(x[10]), .I5(x[11]), .O(n567)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h701F8830CC42A6AA)) n568_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n568)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0CF8FCEFBD9BBBD4)) n569_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n569)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC37C3731808FEE17)) n570_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n570)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h61C19377081F0CEC)) n571_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n571)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n572_lut (
        .I0(n568), .I1(n569), .I2(n570), .I3(n571), .I4(x[6]), .I5(x[10]), .O(n572)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE71113F8444DAD54)) n573_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n573)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF81F094664D2D)) n574_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n574)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h376EEEE77FFFF70C)) n575_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n575)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE3C3C3E8E70F0F80)) n576_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n576)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n577_lut (
        .I0(n573), .I1(n574), .I2(n575), .I3(n576), .I4(x[8]), .I5(x[11]), .O(n577)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4D9C1FC36FA6BE65)) n578_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n578)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2CCE0503D019AA6D)) n579_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n579)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3671E000FFC6CA83)) n580_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n580)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC99C7FAFD7E32FF8)) n581_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[11]), .O(n581)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n582_lut (
        .I0(n578), .I1(n579), .I2(n580), .I3(n581), .I4(x[2]), .I5(x[10]), .O(n582)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6354C70BF35E73CB)) n583_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n583)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1802330F3807A69A)) n584_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n584)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h26813400C03D2541)) n585_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n585)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hDB78F3C000B0CA55)) n586_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n586)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n587_lut (
        .I0(n583), .I1(n584), .I2(n585), .I3(n586), .I4(x[2]), .I5(x[7]), .O(n587)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n588_lut (
        .I0(n572), .I1(n577), .I2(n582), .I3(n587), .I4(x[3]), .I5(x[4]), .O(n588)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFCCF07CB7E4A995)) n589_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n589)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC3C6C00E4A194595)) n590_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n590)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2661E002D33C3F0B)) n591_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n591)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h939C7FFFC98C000F)) n592_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n592)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n593_lut (
        .I0(n589), .I1(n590), .I2(n591), .I3(n592), .I4(x[2]), .I5(x[11]), .O(n593)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE750CF0DF3E37225)) n594_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n594)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h380BC73C73F8A66D)) n595_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n595)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6C810C00000B9556)) n596_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n596)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB3FA3C80003F2FBA)) n597_lut (
        .I0(x[1]), .I1(x[5]), .I2(x[6]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n597)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n598_lut (
        .I0(n594), .I1(n595), .I2(n596), .I3(n597), .I4(x[2]), .I5(x[7]), .O(n598)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC8E0107C462D24AA)) n599_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n599)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0803E7013D4D6296)) n600_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n600)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3C3613310F03CCF0)) n601_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n601)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h9C3CC933E71FFEEF)) n602_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n602)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n603_lut (
        .I0(n599), .I1(n600), .I2(n601), .I3(n602), .I4(x[6]), .I5(x[11]), .O(n603)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3C67E0003CC1966A)) n604_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n604)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h68EEC3FFE0FE262D)) n605_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n605)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6976F3FFFFEF62DB)) n606_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n606)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3C93181FEF3894BD)) n607_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[8]), .I4(x[10]), .I5(x[11]), .O(n607)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n608_lut (
        .I0(n604), .I1(n605), .I2(n606), .I3(n607), .I4(x[6]), .I5(x[7]), .O(n608)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n609_lut (
        .I0(n593), .I1(n598), .I2(n603), .I3(n608), .I4(x[3]), .I5(x[4]), .O(n609)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFF04BF500EA)) n610_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n610)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000030F420057)) n611_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n611)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFE80AB544C243333)) n612_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n612)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5FAA2AFDB3933333)) n613_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n613)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n614_lut (
        .I0(n610), .I1(n611), .I2(n612), .I3(n613), .I4(x[5]), .I5(x[11]), .O(n614)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB4BC2F42FFFFAA05)) n615_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n615)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000803F01F0)) n616_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n616)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCD32CDB33333319C)) n617_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n617)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA801555FD55400AB)) n618_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n618)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n619_lut (
        .I0(n615), .I1(n616), .I2(n617), .I3(n618), .I4(x[10]), .I5(x[11]), .O(n619)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCC9333330AF55000)) n620_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n620)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2CB2CB2C4CB2C34B)) n621_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n621)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000000FFF)) n622_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n622)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h815FA8050FE00FFE)) n623_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[11]), .O(n623)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n624_lut (
        .I0(n620), .I1(n621), .I2(n622), .I3(n623), .I4(x[8]), .I5(x[10]), .O(n624)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h36CB2D34F502AFFF)) n625_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n625)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0FF00FFF000003FF)) n626_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n626)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD2CB2CB224CCD9B3)) n627_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n627)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FA015FEFFFFFFFF)) n628_lut (
        .I0(x[1]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[8]), .O(n628)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n629_lut (
        .I0(n625), .I1(n626), .I2(n627), .I3(n628), .I4(x[10]), .I5(x[11]), .O(n629)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n630_lut (
        .I0(n614), .I1(n619), .I2(n624), .I3(n629), .I4(x[2]), .I5(x[7]), .O(n630)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC13E3CE3E699B3C9)) n631_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n631)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h176878C6C639936C)) n632_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n632)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC1131781EE8800CC)) n633_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n633)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h977EFC7E0177FF73)) n634_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n634)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n635_lut (
        .I0(n631), .I1(n632), .I2(n633), .I3(n634), .I4(x[3]), .I5(x[11]), .O(n635)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h37C800889C339936)) n636_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n636)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC833FFF739339936)) n637_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n637)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h837CE8EC177C1E39)) n638_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n638)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3EC18381ECC17861)) n639_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[11]), .O(n639)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n640_lut (
        .I0(n636), .I1(n637), .I2(n638), .I3(n639), .I4(x[3]), .I5(x[8]), .O(n640)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8CCC6733C00000FF)) n641_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n641)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h33339999FFFF0000)) n642_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n642)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6CCC9999FFFFFFFF)) n643_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n643)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h26649B3301FF0000)) n644_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[6]), .I5(x[11]), .O(n644)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n645_lut (
        .I0(n641), .I1(n642), .I2(n643), .I3(n644), .I4(x[7]), .I5(x[8]), .O(n645)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0080FFFFFFE0FFF8)) n646_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n646)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFF7FFF)) n647_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n647)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB39966999B399966)) n648_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n648)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h99CC26CD993399CE)) n649_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n649)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n650_lut (
        .I0(n646), .I1(n647), .I2(n648), .I3(n649), .I4(x[4]), .I5(x[11]), .O(n650)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n651_lut (
        .I0(n635), .I1(n640), .I2(n645), .I3(n650), .I4(x[5]), .I5(x[10]), .O(n651)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n652_lut (
        .I0(n588), .I1(n609), .I2(n630), .I3(n651), .I4(x[0]), .I5(x[9]), .O(n652)
    );

    wire [10:0] ldtc_tss;
    wire [0:0] ldtc_td;
    assign ldtc_tss[0] = n81;
    assign ldtc_tss[1] = n165;
    assign ldtc_tss[2] = n248;
    assign ldtc_tss[3] = n328;
    assign ldtc_tss[4] = n405;
    assign ldtc_tss[5] = n473;
    assign ldtc_tss[6] = n516;
    assign ldtc_tss[7] = n540;
    assign ldtc_tss[8] = n555;
    assign ldtc_tss[9] = n562;
    assign ldtc_tss[10] = n567;
    assign ldtc_td[0] = n652;
    wire [11:0] ldtc_tss_ext = { { 1{1'b0} }, ldtc_tss } << 1;
    wire [11:0] ldtc_td_ext  = { { 11{1'b0} }, ldtc_td  };
    assign f = ldtc_tss_ext + ldtc_td_ext;
endmodule
