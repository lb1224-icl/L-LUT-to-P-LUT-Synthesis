`timescale 1ns/1ps
module top (input wire [11:0] x, output wire [11:0] f);
    (* KEEP = "TRUE" *) wire n0;
    (* KEEP = "TRUE" *) wire n1;
    (* KEEP = "TRUE" *) wire n2;
    (* KEEP = "TRUE" *) wire n3;
    (* KEEP = "TRUE" *) wire n4;
    (* KEEP = "TRUE" *) wire n5;
    (* KEEP = "TRUE" *) wire n6;
    (* KEEP = "TRUE" *) wire n7;
    (* KEEP = "TRUE" *) wire n8;
    (* KEEP = "TRUE" *) wire n9;
    (* KEEP = "TRUE" *) wire n10;
    (* KEEP = "TRUE" *) wire n11;
    (* KEEP = "TRUE" *) wire n12;
    (* KEEP = "TRUE" *) wire n13;
    (* KEEP = "TRUE" *) wire n14;
    (* KEEP = "TRUE" *) wire n15;
    (* KEEP = "TRUE" *) wire n16;
    (* KEEP = "TRUE" *) wire n17;
    (* KEEP = "TRUE" *) wire n18;
    (* KEEP = "TRUE" *) wire n19;
    (* KEEP = "TRUE" *) wire n20;
    (* KEEP = "TRUE" *) wire n21;
    (* KEEP = "TRUE" *) wire n22;
    (* KEEP = "TRUE" *) wire n23;
    (* KEEP = "TRUE" *) wire n24;
    (* KEEP = "TRUE" *) wire n25;
    (* KEEP = "TRUE" *) wire n26;
    (* KEEP = "TRUE" *) wire n27;
    (* KEEP = "TRUE" *) wire n28;
    (* KEEP = "TRUE" *) wire n29;
    (* KEEP = "TRUE" *) wire n30;
    (* KEEP = "TRUE" *) wire n31;
    (* KEEP = "TRUE" *) wire n32;
    (* KEEP = "TRUE" *) wire n33;
    (* KEEP = "TRUE" *) wire n34;
    (* KEEP = "TRUE" *) wire n35;
    (* KEEP = "TRUE" *) wire n36;
    (* KEEP = "TRUE" *) wire n37;
    (* KEEP = "TRUE" *) wire n38;
    (* KEEP = "TRUE" *) wire n39;
    (* KEEP = "TRUE" *) wire n40;
    (* KEEP = "TRUE" *) wire n41;
    (* KEEP = "TRUE" *) wire n42;
    (* KEEP = "TRUE" *) wire n43;
    (* KEEP = "TRUE" *) wire n44;
    (* KEEP = "TRUE" *) wire n45;
    (* KEEP = "TRUE" *) wire n46;
    (* KEEP = "TRUE" *) wire n47;
    (* KEEP = "TRUE" *) wire n48;
    (* KEEP = "TRUE" *) wire n49;
    (* KEEP = "TRUE" *) wire n50;
    (* KEEP = "TRUE" *) wire n51;
    (* KEEP = "TRUE" *) wire n52;
    (* KEEP = "TRUE" *) wire n53;
    (* KEEP = "TRUE" *) wire n54;
    (* KEEP = "TRUE" *) wire n55;
    (* KEEP = "TRUE" *) wire n56;
    (* KEEP = "TRUE" *) wire n57;
    (* KEEP = "TRUE" *) wire n58;
    (* KEEP = "TRUE" *) wire n59;
    (* KEEP = "TRUE" *) wire n60;
    (* KEEP = "TRUE" *) wire n61;
    (* KEEP = "TRUE" *) wire n62;
    (* KEEP = "TRUE" *) wire n63;
    (* KEEP = "TRUE" *) wire n64;
    (* KEEP = "TRUE" *) wire n65;
    (* KEEP = "TRUE" *) wire n66;
    (* KEEP = "TRUE" *) wire n67;
    (* KEEP = "TRUE" *) wire n68;
    (* KEEP = "TRUE" *) wire n69;
    (* KEEP = "TRUE" *) wire n70;
    (* KEEP = "TRUE" *) wire n71;
    (* KEEP = "TRUE" *) wire n72;
    (* KEEP = "TRUE" *) wire n73;
    (* KEEP = "TRUE" *) wire n74;
    (* KEEP = "TRUE" *) wire n75;
    (* KEEP = "TRUE" *) wire n76;
    (* KEEP = "TRUE" *) wire n77;
    (* KEEP = "TRUE" *) wire n78;
    (* KEEP = "TRUE" *) wire n79;
    (* KEEP = "TRUE" *) wire n80;
    (* KEEP = "TRUE" *) wire n81;
    (* KEEP = "TRUE" *) wire n82;
    (* KEEP = "TRUE" *) wire n83;
    (* KEEP = "TRUE" *) wire n84;
    (* KEEP = "TRUE" *) wire n85;
    (* KEEP = "TRUE" *) wire n86;
    (* KEEP = "TRUE" *) wire n87;
    (* KEEP = "TRUE" *) wire n88;
    (* KEEP = "TRUE" *) wire n89;
    (* KEEP = "TRUE" *) wire n90;
    (* KEEP = "TRUE" *) wire n91;
    (* KEEP = "TRUE" *) wire n92;
    (* KEEP = "TRUE" *) wire n93;
    (* KEEP = "TRUE" *) wire n94;
    (* KEEP = "TRUE" *) wire n95;
    (* KEEP = "TRUE" *) wire n96;
    (* KEEP = "TRUE" *) wire n97;
    (* KEEP = "TRUE" *) wire n98;
    (* KEEP = "TRUE" *) wire n99;
    (* KEEP = "TRUE" *) wire n100;
    (* KEEP = "TRUE" *) wire n101;
    (* KEEP = "TRUE" *) wire n102;
    (* KEEP = "TRUE" *) wire n103;
    (* KEEP = "TRUE" *) wire n104;
    (* KEEP = "TRUE" *) wire n105;
    (* KEEP = "TRUE" *) wire n106;
    (* KEEP = "TRUE" *) wire n107;
    (* KEEP = "TRUE" *) wire n108;
    (* KEEP = "TRUE" *) wire n109;
    (* KEEP = "TRUE" *) wire n110;
    (* KEEP = "TRUE" *) wire n111;
    (* KEEP = "TRUE" *) wire n112;
    (* KEEP = "TRUE" *) wire n113;
    (* KEEP = "TRUE" *) wire n114;
    (* KEEP = "TRUE" *) wire n115;
    (* KEEP = "TRUE" *) wire n116;
    (* KEEP = "TRUE" *) wire n117;
    (* KEEP = "TRUE" *) wire n118;
    (* KEEP = "TRUE" *) wire n119;
    (* KEEP = "TRUE" *) wire n120;
    (* KEEP = "TRUE" *) wire n121;
    (* KEEP = "TRUE" *) wire n122;
    (* KEEP = "TRUE" *) wire n123;
    (* KEEP = "TRUE" *) wire n124;
    (* KEEP = "TRUE" *) wire n125;
    (* KEEP = "TRUE" *) wire n126;
    (* KEEP = "TRUE" *) wire n127;
    (* KEEP = "TRUE" *) wire n128;
    (* KEEP = "TRUE" *) wire n129;
    (* KEEP = "TRUE" *) wire n130;
    (* KEEP = "TRUE" *) wire n131;
    (* KEEP = "TRUE" *) wire n132;
    (* KEEP = "TRUE" *) wire n133;
    (* KEEP = "TRUE" *) wire n134;
    (* KEEP = "TRUE" *) wire n135;
    (* KEEP = "TRUE" *) wire n136;
    (* KEEP = "TRUE" *) wire n137;
    (* KEEP = "TRUE" *) wire n138;
    (* KEEP = "TRUE" *) wire n139;
    (* KEEP = "TRUE" *) wire n140;
    (* KEEP = "TRUE" *) wire n141;
    (* KEEP = "TRUE" *) wire n142;
    (* KEEP = "TRUE" *) wire n143;
    (* KEEP = "TRUE" *) wire n144;
    (* KEEP = "TRUE" *) wire n145;
    (* KEEP = "TRUE" *) wire n146;
    (* KEEP = "TRUE" *) wire n147;
    (* KEEP = "TRUE" *) wire n148;
    (* KEEP = "TRUE" *) wire n149;
    (* KEEP = "TRUE" *) wire n150;
    (* KEEP = "TRUE" *) wire n151;
    (* KEEP = "TRUE" *) wire n152;
    (* KEEP = "TRUE" *) wire n153;
    (* KEEP = "TRUE" *) wire n154;
    (* KEEP = "TRUE" *) wire n155;
    (* KEEP = "TRUE" *) wire n156;
    (* KEEP = "TRUE" *) wire n157;
    (* KEEP = "TRUE" *) wire n158;
    (* KEEP = "TRUE" *) wire n159;
    (* KEEP = "TRUE" *) wire n160;
    (* KEEP = "TRUE" *) wire n161;
    (* KEEP = "TRUE" *) wire n162;
    (* KEEP = "TRUE" *) wire n163;
    (* KEEP = "TRUE" *) wire n164;
    (* KEEP = "TRUE" *) wire n165;
    (* KEEP = "TRUE" *) wire n166;
    (* KEEP = "TRUE" *) wire n167;
    (* KEEP = "TRUE" *) wire n168;
    (* KEEP = "TRUE" *) wire n169;
    (* KEEP = "TRUE" *) wire n170;
    (* KEEP = "TRUE" *) wire n171;
    (* KEEP = "TRUE" *) wire n172;
    (* KEEP = "TRUE" *) wire n173;
    (* KEEP = "TRUE" *) wire n174;
    (* KEEP = "TRUE" *) wire n175;
    (* KEEP = "TRUE" *) wire n176;
    (* KEEP = "TRUE" *) wire n177;
    (* KEEP = "TRUE" *) wire n178;
    (* KEEP = "TRUE" *) wire n179;
    (* KEEP = "TRUE" *) wire n180;
    (* KEEP = "TRUE" *) wire n181;
    (* KEEP = "TRUE" *) wire n182;
    (* KEEP = "TRUE" *) wire n183;
    (* KEEP = "TRUE" *) wire n184;
    (* KEEP = "TRUE" *) wire n185;
    (* KEEP = "TRUE" *) wire n186;
    (* KEEP = "TRUE" *) wire n187;
    (* KEEP = "TRUE" *) wire n188;
    (* KEEP = "TRUE" *) wire n189;
    (* KEEP = "TRUE" *) wire n190;
    (* KEEP = "TRUE" *) wire n191;
    (* KEEP = "TRUE" *) wire n192;
    (* KEEP = "TRUE" *) wire n193;
    (* KEEP = "TRUE" *) wire n194;
    (* KEEP = "TRUE" *) wire n195;
    (* KEEP = "TRUE" *) wire n196;
    (* KEEP = "TRUE" *) wire n197;
    (* KEEP = "TRUE" *) wire n198;
    (* KEEP = "TRUE" *) wire n199;
    (* KEEP = "TRUE" *) wire n200;
    (* KEEP = "TRUE" *) wire n201;
    (* KEEP = "TRUE" *) wire n202;
    (* KEEP = "TRUE" *) wire n203;
    (* KEEP = "TRUE" *) wire n204;
    (* KEEP = "TRUE" *) wire n205;
    (* KEEP = "TRUE" *) wire n206;
    (* KEEP = "TRUE" *) wire n207;
    (* KEEP = "TRUE" *) wire n208;
    (* KEEP = "TRUE" *) wire n209;
    (* KEEP = "TRUE" *) wire n210;
    (* KEEP = "TRUE" *) wire n211;
    (* KEEP = "TRUE" *) wire n212;
    (* KEEP = "TRUE" *) wire n213;
    (* KEEP = "TRUE" *) wire n214;
    (* KEEP = "TRUE" *) wire n215;
    (* KEEP = "TRUE" *) wire n216;
    (* KEEP = "TRUE" *) wire n217;
    (* KEEP = "TRUE" *) wire n218;
    (* KEEP = "TRUE" *) wire n219;
    (* KEEP = "TRUE" *) wire n220;
    (* KEEP = "TRUE" *) wire n221;
    (* KEEP = "TRUE" *) wire n222;
    (* KEEP = "TRUE" *) wire n223;
    (* KEEP = "TRUE" *) wire n224;
    (* KEEP = "TRUE" *) wire n225;
    (* KEEP = "TRUE" *) wire n226;
    (* KEEP = "TRUE" *) wire n227;
    (* KEEP = "TRUE" *) wire n228;
    (* KEEP = "TRUE" *) wire n229;
    (* KEEP = "TRUE" *) wire n230;
    (* KEEP = "TRUE" *) wire n231;
    (* KEEP = "TRUE" *) wire n232;
    (* KEEP = "TRUE" *) wire n233;
    (* KEEP = "TRUE" *) wire n234;
    (* KEEP = "TRUE" *) wire n235;
    (* KEEP = "TRUE" *) wire n236;
    (* KEEP = "TRUE" *) wire n237;
    (* KEEP = "TRUE" *) wire n238;
    (* KEEP = "TRUE" *) wire n239;
    (* KEEP = "TRUE" *) wire n240;
    (* KEEP = "TRUE" *) wire n241;
    (* KEEP = "TRUE" *) wire n242;
    (* KEEP = "TRUE" *) wire n243;
    (* KEEP = "TRUE" *) wire n244;
    (* KEEP = "TRUE" *) wire n245;
    (* KEEP = "TRUE" *) wire n246;
    (* KEEP = "TRUE" *) wire n247;
    (* KEEP = "TRUE" *) wire n248;
    (* KEEP = "TRUE" *) wire n249;
    (* KEEP = "TRUE" *) wire n250;
    (* KEEP = "TRUE" *) wire n251;
    (* KEEP = "TRUE" *) wire n252;
    (* KEEP = "TRUE" *) wire n253;
    (* KEEP = "TRUE" *) wire n254;
    (* KEEP = "TRUE" *) wire n255;
    (* KEEP = "TRUE" *) wire n256;
    (* KEEP = "TRUE" *) wire n257;
    (* KEEP = "TRUE" *) wire n258;
    (* KEEP = "TRUE" *) wire n259;
    (* KEEP = "TRUE" *) wire n260;
    (* KEEP = "TRUE" *) wire n261;
    (* KEEP = "TRUE" *) wire n262;
    (* KEEP = "TRUE" *) wire n263;
    (* KEEP = "TRUE" *) wire n264;
    (* KEEP = "TRUE" *) wire n265;
    (* KEEP = "TRUE" *) wire n266;
    (* KEEP = "TRUE" *) wire n267;
    (* KEEP = "TRUE" *) wire n268;
    (* KEEP = "TRUE" *) wire n269;
    (* KEEP = "TRUE" *) wire n270;
    (* KEEP = "TRUE" *) wire n271;
    (* KEEP = "TRUE" *) wire n272;
    (* KEEP = "TRUE" *) wire n273;
    (* KEEP = "TRUE" *) wire n274;
    (* KEEP = "TRUE" *) wire n275;
    (* KEEP = "TRUE" *) wire n276;
    (* KEEP = "TRUE" *) wire n277;
    (* KEEP = "TRUE" *) wire n278;
    (* KEEP = "TRUE" *) wire n279;
    (* KEEP = "TRUE" *) wire n280;
    (* KEEP = "TRUE" *) wire n281;
    (* KEEP = "TRUE" *) wire n282;
    (* KEEP = "TRUE" *) wire n283;
    (* KEEP = "TRUE" *) wire n284;
    (* KEEP = "TRUE" *) wire n285;
    (* KEEP = "TRUE" *) wire n286;
    (* KEEP = "TRUE" *) wire n287;
    (* KEEP = "TRUE" *) wire n288;
    (* KEEP = "TRUE" *) wire n289;
    (* KEEP = "TRUE" *) wire n290;
    (* KEEP = "TRUE" *) wire n291;
    (* KEEP = "TRUE" *) wire n292;
    (* KEEP = "TRUE" *) wire n293;
    (* KEEP = "TRUE" *) wire n294;
    (* KEEP = "TRUE" *) wire n295;
    (* KEEP = "TRUE" *) wire n296;
    (* KEEP = "TRUE" *) wire n297;
    (* KEEP = "TRUE" *) wire n298;
    (* KEEP = "TRUE" *) wire n299;
    (* KEEP = "TRUE" *) wire n300;
    (* KEEP = "TRUE" *) wire n301;
    (* KEEP = "TRUE" *) wire n302;
    (* KEEP = "TRUE" *) wire n303;
    (* KEEP = "TRUE" *) wire n304;
    (* KEEP = "TRUE" *) wire n305;
    (* KEEP = "TRUE" *) wire n306;
    (* KEEP = "TRUE" *) wire n307;
    (* KEEP = "TRUE" *) wire n308;
    (* KEEP = "TRUE" *) wire n309;
    (* KEEP = "TRUE" *) wire n310;
    (* KEEP = "TRUE" *) wire n311;
    (* KEEP = "TRUE" *) wire n312;
    (* KEEP = "TRUE" *) wire n313;
    (* KEEP = "TRUE" *) wire n314;
    (* KEEP = "TRUE" *) wire n315;
    (* KEEP = "TRUE" *) wire n316;
    (* KEEP = "TRUE" *) wire n317;
    (* KEEP = "TRUE" *) wire n318;
    (* KEEP = "TRUE" *) wire n319;
    (* KEEP = "TRUE" *) wire n320;
    (* KEEP = "TRUE" *) wire n321;
    (* KEEP = "TRUE" *) wire n322;
    (* KEEP = "TRUE" *) wire n323;
    (* KEEP = "TRUE" *) wire n324;
    (* KEEP = "TRUE" *) wire n325;
    (* KEEP = "TRUE" *) wire n326;
    (* KEEP = "TRUE" *) wire n327;
    (* KEEP = "TRUE" *) wire n328;
    (* KEEP = "TRUE" *) wire n329;
    (* KEEP = "TRUE" *) wire n330;
    (* KEEP = "TRUE" *) wire n331;
    (* KEEP = "TRUE" *) wire n332;
    (* KEEP = "TRUE" *) wire n333;
    (* KEEP = "TRUE" *) wire n334;
    (* KEEP = "TRUE" *) wire n335;
    (* KEEP = "TRUE" *) wire n336;
    (* KEEP = "TRUE" *) wire n337;
    (* KEEP = "TRUE" *) wire n338;
    (* KEEP = "TRUE" *) wire n339;
    (* KEEP = "TRUE" *) wire n340;
    (* KEEP = "TRUE" *) wire n341;
    (* KEEP = "TRUE" *) wire n342;
    (* KEEP = "TRUE" *) wire n343;
    (* KEEP = "TRUE" *) wire n344;
    (* KEEP = "TRUE" *) wire n345;
    (* KEEP = "TRUE" *) wire n346;
    (* KEEP = "TRUE" *) wire n347;
    (* KEEP = "TRUE" *) wire n348;
    (* KEEP = "TRUE" *) wire n349;
    (* KEEP = "TRUE" *) wire n350;
    (* KEEP = "TRUE" *) wire n351;
    (* KEEP = "TRUE" *) wire n352;
    (* KEEP = "TRUE" *) wire n353;
    (* KEEP = "TRUE" *) wire n354;
    (* KEEP = "TRUE" *) wire n355;
    (* KEEP = "TRUE" *) wire n356;
    (* KEEP = "TRUE" *) wire n357;
    (* KEEP = "TRUE" *) wire n358;
    (* KEEP = "TRUE" *) wire n359;
    (* KEEP = "TRUE" *) wire n360;
    (* KEEP = "TRUE" *) wire n361;
    (* KEEP = "TRUE" *) wire n362;
    (* KEEP = "TRUE" *) wire n363;
    (* KEEP = "TRUE" *) wire n364;
    (* KEEP = "TRUE" *) wire n365;
    (* KEEP = "TRUE" *) wire n366;
    (* KEEP = "TRUE" *) wire n367;
    (* KEEP = "TRUE" *) wire n368;
    (* KEEP = "TRUE" *) wire n369;
    (* KEEP = "TRUE" *) wire n370;
    (* KEEP = "TRUE" *) wire n371;
    (* KEEP = "TRUE" *) wire n372;
    (* KEEP = "TRUE" *) wire n373;
    (* KEEP = "TRUE" *) wire n374;
    (* KEEP = "TRUE" *) wire n375;
    (* KEEP = "TRUE" *) wire n376;
    (* KEEP = "TRUE" *) wire n377;
    (* KEEP = "TRUE" *) wire n378;
    (* KEEP = "TRUE" *) wire n379;
    (* KEEP = "TRUE" *) wire n380;
    (* KEEP = "TRUE" *) wire n381;
    (* KEEP = "TRUE" *) wire n382;
    (* KEEP = "TRUE" *) wire n383;
    (* KEEP = "TRUE" *) wire n384;
    (* KEEP = "TRUE" *) wire n385;
    (* KEEP = "TRUE" *) wire n386;
    (* KEEP = "TRUE" *) wire n387;
    (* KEEP = "TRUE" *) wire n388;
    (* KEEP = "TRUE" *) wire n389;
    (* KEEP = "TRUE" *) wire n390;
    (* KEEP = "TRUE" *) wire n391;
    (* KEEP = "TRUE" *) wire n392;
    (* KEEP = "TRUE" *) wire n393;
    (* KEEP = "TRUE" *) wire n394;
    (* KEEP = "TRUE" *) wire n395;
    (* KEEP = "TRUE" *) wire n396;
    (* KEEP = "TRUE" *) wire n397;
    (* KEEP = "TRUE" *) wire n398;
    (* KEEP = "TRUE" *) wire n399;
    (* KEEP = "TRUE" *) wire n400;
    (* KEEP = "TRUE" *) wire n401;
    (* KEEP = "TRUE" *) wire n402;
    (* KEEP = "TRUE" *) wire n403;
    (* KEEP = "TRUE" *) wire n404;
    (* KEEP = "TRUE" *) wire n405;
    (* KEEP = "TRUE" *) wire n406;
    (* KEEP = "TRUE" *) wire n407;
    (* KEEP = "TRUE" *) wire n408;
    (* KEEP = "TRUE" *) wire n409;
    (* KEEP = "TRUE" *) wire n410;
    (* KEEP = "TRUE" *) wire n411;
    (* KEEP = "TRUE" *) wire n412;
    (* KEEP = "TRUE" *) wire n413;
    (* KEEP = "TRUE" *) wire n414;
    (* KEEP = "TRUE" *) wire n415;
    (* KEEP = "TRUE" *) wire n416;
    (* KEEP = "TRUE" *) wire n417;
    (* KEEP = "TRUE" *) wire n418;
    (* KEEP = "TRUE" *) wire n419;
    (* KEEP = "TRUE" *) wire n420;
    (* KEEP = "TRUE" *) wire n421;
    (* KEEP = "TRUE" *) wire n422;
    (* KEEP = "TRUE" *) wire n423;
    (* KEEP = "TRUE" *) wire n424;
    (* KEEP = "TRUE" *) wire n425;
    (* KEEP = "TRUE" *) wire n426;
    (* KEEP = "TRUE" *) wire n427;
    (* KEEP = "TRUE" *) wire n428;
    (* KEEP = "TRUE" *) wire n429;
    (* KEEP = "TRUE" *) wire n430;
    (* KEEP = "TRUE" *) wire n431;
    (* KEEP = "TRUE" *) wire n432;
    (* KEEP = "TRUE" *) wire n433;
    (* KEEP = "TRUE" *) wire n434;
    (* KEEP = "TRUE" *) wire n435;
    (* KEEP = "TRUE" *) wire n436;
    (* KEEP = "TRUE" *) wire n437;
    (* KEEP = "TRUE" *) wire n438;
    (* KEEP = "TRUE" *) wire n439;
    (* KEEP = "TRUE" *) wire n440;
    (* KEEP = "TRUE" *) wire n441;
    (* KEEP = "TRUE" *) wire n442;
    (* KEEP = "TRUE" *) wire n443;
    (* KEEP = "TRUE" *) wire n444;
    (* KEEP = "TRUE" *) wire n445;
    (* KEEP = "TRUE" *) wire n446;
    (* KEEP = "TRUE" *) wire n447;
    (* KEEP = "TRUE" *) wire n448;
    (* KEEP = "TRUE" *) wire n449;
    (* KEEP = "TRUE" *) wire n450;
    (* KEEP = "TRUE" *) wire n451;
    (* KEEP = "TRUE" *) wire n452;
    (* KEEP = "TRUE" *) wire n453;
    (* KEEP = "TRUE" *) wire n454;
    (* KEEP = "TRUE" *) wire n455;
    (* KEEP = "TRUE" *) wire n456;
    (* KEEP = "TRUE" *) wire n457;
    (* KEEP = "TRUE" *) wire n458;
    (* KEEP = "TRUE" *) wire n459;
    (* KEEP = "TRUE" *) wire n460;
    (* KEEP = "TRUE" *) wire n461;
    (* KEEP = "TRUE" *) wire n462;
    (* KEEP = "TRUE" *) wire n463;
    (* KEEP = "TRUE" *) wire n464;
    (* KEEP = "TRUE" *) wire n465;
    (* KEEP = "TRUE" *) wire n466;
    (* KEEP = "TRUE" *) wire n467;
    (* KEEP = "TRUE" *) wire n468;
    (* KEEP = "TRUE" *) wire n469;
    (* KEEP = "TRUE" *) wire n470;
    (* KEEP = "TRUE" *) wire n471;
    (* KEEP = "TRUE" *) wire n472;
    (* KEEP = "TRUE" *) wire n473;
    (* KEEP = "TRUE" *) wire n474;
    (* KEEP = "TRUE" *) wire n475;
    (* KEEP = "TRUE" *) wire n476;
    (* KEEP = "TRUE" *) wire n477;
    (* KEEP = "TRUE" *) wire n478;
    (* KEEP = "TRUE" *) wire n479;
    (* KEEP = "TRUE" *) wire n480;
    (* KEEP = "TRUE" *) wire n481;
    (* KEEP = "TRUE" *) wire n482;
    (* KEEP = "TRUE" *) wire n483;
    (* KEEP = "TRUE" *) wire n484;
    (* KEEP = "TRUE" *) wire n485;
    (* KEEP = "TRUE" *) wire n486;
    (* KEEP = "TRUE" *) wire n487;
    (* KEEP = "TRUE" *) wire n488;
    (* KEEP = "TRUE" *) wire n489;
    (* KEEP = "TRUE" *) wire n490;
    (* KEEP = "TRUE" *) wire n491;
    (* KEEP = "TRUE" *) wire n492;
    (* KEEP = "TRUE" *) wire n493;
    (* KEEP = "TRUE" *) wire n494;
    (* KEEP = "TRUE" *) wire n495;
    (* KEEP = "TRUE" *) wire n496;
    (* KEEP = "TRUE" *) wire n497;
    (* KEEP = "TRUE" *) wire n498;
    (* KEEP = "TRUE" *) wire n499;
    (* KEEP = "TRUE" *) wire n500;
    (* KEEP = "TRUE" *) wire n501;
    (* KEEP = "TRUE" *) wire n502;
    (* KEEP = "TRUE" *) wire n503;
    (* KEEP = "TRUE" *) wire n504;
    (* KEEP = "TRUE" *) wire n505;
    (* KEEP = "TRUE" *) wire n506;
    (* KEEP = "TRUE" *) wire n507;
    (* KEEP = "TRUE" *) wire n508;
    (* KEEP = "TRUE" *) wire n509;
    (* KEEP = "TRUE" *) wire n510;
    (* KEEP = "TRUE" *) wire n511;
    (* KEEP = "TRUE" *) wire n512;
    (* KEEP = "TRUE" *) wire n513;
    (* KEEP = "TRUE" *) wire n514;
    (* KEEP = "TRUE" *) wire n515;
    (* KEEP = "TRUE" *) wire n516;
    (* KEEP = "TRUE" *) wire n517;
    (* KEEP = "TRUE" *) wire n518;
    (* KEEP = "TRUE" *) wire n519;
    (* KEEP = "TRUE" *) wire n520;
    (* KEEP = "TRUE" *) wire n521;
    (* KEEP = "TRUE" *) wire n522;
    (* KEEP = "TRUE" *) wire n523;

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h33FF68FF1FF15A5A)) n0_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n0)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA6B4A5426C8155A5)) n1_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n1)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h95AD6655A55B22A5)) n2_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n2)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD2B5FFFFEE6CE396)) n3_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n3)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n4_lut (
        .I0(n0), .I1(n1), .I2(n2), .I3(n3), .I4(x[7]), .I5(x[8]), .O(n4)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h30E04017AC62530C)) n5_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n5)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCF9847E3517296FB)) n6_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n6)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h33F53A195D23377E)) n7_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n7)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCC25396902639A89)) n8_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n8)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n9_lut (
        .I0(n5), .I1(n6), .I2(n7), .I3(n8), .I4(x[1]), .I5(x[6]), .O(n9)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA04501F825605B00)) n10_lut (
        .I0(x[2]), .I1(x[6]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n10)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5D950A081E9864FF)) n11_lut (
        .I0(x[2]), .I1(x[6]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n11)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h73A6FA48C0675E3F)) n12_lut (
        .I0(x[2]), .I1(x[6]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n12)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEC5A7D98E5E329C0)) n13_lut (
        .I0(x[2]), .I1(x[6]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n13)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n14_lut (
        .I0(n10), .I1(n11), .I2(n12), .I3(n13), .I4(x[1]), .I5(x[4]), .O(n14)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD39E6CFFEFFE5A96)) n15_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n15)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5A99A55B44CC6A52)) n16_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n16)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4A55036C945A4BDB)) n17_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n17)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA5A50EF0FF3CEE99)) n18_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n18)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n19_lut (
        .I0(n15), .I1(n16), .I2(n17), .I3(n18), .I4(x[7]), .I5(x[8]), .O(n19)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n20_lut (
        .I0(n4), .I1(n9), .I2(n14), .I3(n19), .I4(x[3]), .I5(x[5]), .O(n20)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h64AA8EFF3CBDA595)) n21_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n21)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h86AD37003652AD42)) n22_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n22)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0E962B30CED5AADB)) n23_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n23)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFBB6DFEF1355AA6)) n24_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n24)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n25_lut (
        .I0(n21), .I1(n22), .I2(n23), .I3(n24), .I4(x[4]), .I5(x[6]), .O(n25)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1692610CC0038CCC)) n26_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n26)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h065597D31FFC3333)) n27_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n27)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF46AEB0359584C1D)) n28_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n28)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF03594FCA2680C0C)) n29_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n29)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n30_lut (
        .I0(n26), .I1(n27), .I2(n28), .I3(n29), .I4(x[1]), .I5(x[9]), .O(n30)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h303016453F29AC0F)) n31_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n31)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB8321A9AC0D7562F)) n32_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n32)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCCCC3FF8CBE9AA60)) n33_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n33)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3331C00330864968)) n34_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n34)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n35_lut (
        .I0(n31), .I1(n32), .I2(n33), .I3(n34), .I4(x[1]), .I5(x[9]), .O(n35)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h655AAC8F7FB6DDFF)) n36_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n36)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hDB55AB730CD46970)) n37_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n37)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h42B54A6C00ECB561)) n38_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n38)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA9A5BD3CFF715526)) n39_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n39)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n40_lut (
        .I0(n36), .I1(n37), .I2(n38), .I3(n39), .I4(x[4]), .I5(x[6]), .O(n40)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n41_lut (
        .I0(n25), .I1(n30), .I2(n35), .I3(n40), .I4(x[3]), .I5(x[10]), .O(n41)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCC009700E00EA5A4)) n42_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n42)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n43_lut (
        .I0(n42), .I1(~(n1)), .I2(~(n2)), .I3(~(n3)), .I4(x[7]), .I5(x[8]), .O(n43)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n44_lut (
        .I0(~(n5)), .I1(~(n6)), .I2(~(n7)), .I3(~(n8)), .I4(x[1]), .I5(x[6]), .O(n44)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n45_lut (
        .I0(~(n10)), .I1(~(n11)), .I2(~(n12)), .I3(~(n13)), .I4(x[1]), .I5(x[4]), .O(n45)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n46_lut (
        .I0(~(n15)), .I1(~(n16)), .I2(~(n17)), .I3(~(n18)), .I4(x[7]), .I5(x[8]), .O(n46)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n47_lut (
        .I0(n43), .I1(n44), .I2(n45), .I3(n46), .I4(x[3]), .I5(x[5]), .O(n47)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n48_lut (
        .I0(~(n21)), .I1(~(n22)), .I2(~(n23)), .I3(~(n24)), .I4(x[4]), .I5(x[6]), .O(n48)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n49_lut (
        .I0(~(n26)), .I1(~(n27)), .I2(~(n28)), .I3(~(n29)), .I4(x[1]), .I5(x[9]), .O(n49)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n50_lut (
        .I0(~(n31)), .I1(~(n32)), .I2(~(n33)), .I3(~(n34)), .I4(x[1]), .I5(x[9]), .O(n50)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n51_lut (
        .I0(~(n36)), .I1(~(n37)), .I2(~(n38)), .I3(~(n39)), .I4(x[4]), .I5(x[6]), .O(n51)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n52_lut (
        .I0(n48), .I1(n49), .I2(n50), .I3(n51), .I4(x[3]), .I5(x[10]), .O(n52)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n53_lut (
        .I0(n20), .I1(n41), .I2(n47), .I3(n52), .I4(x[0]), .I5(x[11]), .O(n53)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h9E7FCEFFBDF169BC)) n54_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n54)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h898833CF2BF56634)) n55_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n55)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD3635FCC00D26A69)) n56_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n56)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hD6665FDFFFC11E73)) n57_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n57)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n58_lut (
        .I0(n54), .I1(n55), .I2(n56), .I3(n57), .I4(x[6]), .I5(x[8]), .O(n58)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1AD56803F33C5986)) n59_lut (
        .I0(x[0]), .I1(x[5]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n59)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h656161A3FC668679)) n60_lut (
        .I0(x[0]), .I1(x[5]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n60)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3A7F7CFCD3C91AA6)) n61_lut (
        .I0(x[0]), .I1(x[5]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n61)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h45853810C0999D59)) n62_lut (
        .I0(x[0]), .I1(x[5]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n62)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n63_lut (
        .I0(n59), .I1(n60), .I2(n61), .I3(n62), .I4(x[2]), .I5(x[6]), .O(n63)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0D363EF8EC96C66)) n64_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n64)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F0D33C0E698C699)) n65_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n65)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h99666780003330DA)) n66_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n66)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6666968EF03CDB05)) n67_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n67)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n68_lut (
        .I0(n64), .I1(n65), .I2(n66), .I3(n67), .I4(x[5]), .I5(x[9]), .O(n68)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h542B6E3F79936666)) n69_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n69)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hAF52933F5179869D)) n70_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n70)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h99666E7ACFE9CDFF)) n71_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n71)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h66261815FCC94445)) n72_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n72)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n73_lut (
        .I0(n69), .I1(n70), .I2(n71), .I3(n72), .I4(x[5]), .I5(x[9]), .O(n73)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n74_lut (
        .I0(n58), .I1(n63), .I2(n68), .I3(n73), .I4(x[3]), .I5(x[4]), .O(n74)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7861667199996499)) n75_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n75)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3C38CCD32B50055F)) n76_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n76)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hBF50CB3431C7FFFF)) n77_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n77)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h9366CC669E7917A0)) n78_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[8]), .O(n78)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n79_lut (
        .I0(n75), .I1(n76), .I2(n77), .I3(n78), .I4(x[9]), .I5(x[10]), .O(n79)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5434222300180416)) n80_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n80)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEA9224B13F78ABE9)) n81_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n81)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h156B2D4CB0FAFD16)) n82_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n82)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6A9D0B3CFF8A56F8)) n83_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n83)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n84_lut (
        .I0(n80), .I1(n81), .I2(n82), .I3(n83), .I4(x[2]), .I5(x[3]), .O(n84)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2DBF0A5D36E0D6A9)) n85_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n85)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5A94805D36A309A2)) n86_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n86)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h69600D54C4102C2B)) n87_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n87)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hDA9ACF50C653B6A6)) n88_lut (
        .I0(x[2]), .I1(x[4]), .I2(x[7]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n88)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n89_lut (
        .I0(n85), .I1(n86), .I2(n87), .I3(n88), .I4(x[0]), .I5(x[3]), .O(n89)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h34CBAF5499999366)) n90_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n90)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFF3CEA05EE79E)) n91_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n91)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6739E1A7CD930E1E)) n92_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n92)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6C99666C57FA2F42)) n93_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[7]), .I5(x[9]), .O(n93)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n94_lut (
        .I0(n90), .I1(n91), .I2(n92), .I3(n93), .I4(x[8]), .I5(x[10]), .O(n94)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n95_lut (
        .I0(n79), .I1(n84), .I2(n89), .I3(n94), .I4(x[5]), .I5(x[6]), .O(n95)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h61803100420E9642)) n96_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n96)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n97_lut (
        .I0(n96), .I1(~(n55)), .I2(~(n56)), .I3(~(n57)), .I4(x[6]), .I5(x[8]), .O(n97)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n98_lut (
        .I0(~(n59)), .I1(~(n60)), .I2(~(n61)), .I3(~(n62)), .I4(x[2]), .I5(x[6]), .O(n98)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n99_lut (
        .I0(~(n64)), .I1(~(n65)), .I2(~(n66)), .I3(~(n67)), .I4(x[5]), .I5(x[9]), .O(n99)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n100_lut (
        .I0(~(n69)), .I1(~(n70)), .I2(~(n71)), .I3(~(n72)), .I4(x[5]), .I5(x[9]), .O(n100)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n101_lut (
        .I0(n97), .I1(n98), .I2(n99), .I3(n100), .I4(x[3]), .I5(x[4]), .O(n101)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n102_lut (
        .I0(~(n75)), .I1(~(n76)), .I2(~(n77)), .I3(~(n78)), .I4(x[9]), .I5(x[10]), .O(n102)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n103_lut (
        .I0(~(n80)), .I1(~(n81)), .I2(~(n82)), .I3(~(n83)), .I4(x[2]), .I5(x[3]), .O(n103)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n104_lut (
        .I0(~(n85)), .I1(~(n86)), .I2(~(n87)), .I3(~(n88)), .I4(x[0]), .I5(x[3]), .O(n104)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n105_lut (
        .I0(~(n90)), .I1(~(n91)), .I2(~(n92)), .I3(~(n93)), .I4(x[8]), .I5(x[10]), .O(n105)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n106_lut (
        .I0(n102), .I1(n103), .I2(n104), .I3(n105), .I4(x[5]), .I5(x[6]), .O(n106)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n107_lut (
        .I0(n74), .I1(n95), .I2(n101), .I3(n106), .I4(x[1]), .I5(x[11]), .O(n107)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hABC03C8F205E05F0)) n108_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n108)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFD3C3CCF3C07B21E)) n109_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n109)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hAAC7333FCEF7BF78)) n110_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n110)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7F33D19FCFC0C407)) n111_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n111)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n112_lut (
        .I0(n108), .I1(n109), .I2(n110), .I3(n111), .I4(x[1]), .I5(x[5]), .O(n112)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3463CC3FCB42A05F)) n113_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n113)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB330CC3F2C2F7E81)) n114_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n114)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h555533383F47FD7F)) n115_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n115)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA002938E3C01D001)) n116_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n116)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n117_lut (
        .I0(n113), .I1(n114), .I2(n115), .I3(n116), .I4(x[1]), .I5(x[9]), .O(n117)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7F70008118C88C89)) n118_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n118)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3FF3010FC7338CC8)) n119_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n119)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC9373C3EF0FFF37E)) n120_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n120)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE81331E8FF0018C0)) n121_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n121)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n122_lut (
        .I0(n118), .I1(n119), .I2(n120), .I3(n121), .I4(x[4]), .I5(x[9]), .O(n122)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFDFBF48E66FFFF)) n123_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n123)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h07D0FFF0E3335015)) n124_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n124)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7F800BCBFE33C334)) n125_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n125)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h81FEBD2CFF33F332)) n126_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n126)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n127_lut (
        .I0(n123), .I1(n124), .I2(n125), .I3(n126), .I4(x[1]), .I5(x[9]), .O(n127)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n128_lut (
        .I0(n112), .I1(n117), .I2(n122), .I3(n127), .I4(x[3]), .I5(x[7]), .O(n128)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h70F3EC801133C893)) n129_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n129)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F0FFFFFE1C3CE73)) n130_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n130)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8E38F83F8FF0FFFF)) n131_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n131)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h37EC88CC08CFF07F)) n132_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[7]), .I5(x[9]), .O(n132)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n133_lut (
        .I0(n129), .I1(n130), .I2(n131), .I3(n132), .I4(x[8]), .I5(x[10]), .O(n133)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3EC71EFF17E8EC3E)) n134_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n134)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h6831F00FECECEE36)) n135_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n135)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h81730E30F3008818)) n136_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n136)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC973088E0C007778)) n137_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n137)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n138_lut (
        .I0(n134), .I1(n135), .I2(n136), .I3(n137), .I4(x[4]), .I5(x[8]), .O(n138)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF00F008EF3E8117E)) n139_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n139)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF0F8F0C38833136)) n140_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n140)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h83C8611180000000)) n141_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n141)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC1CCE3EEC83FC0FF)) n142_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[7]), .I4(x[8]), .I5(x[9]), .O(n142)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n143_lut (
        .I0(n139), .I1(n140), .I2(n141), .I3(n142), .I4(x[4]), .I5(x[10]), .O(n143)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F3018CEE38EC891)) n144_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n144)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF1FC117E1CEEE)) n145_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n145)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h33373878F1C7F0F0)) n146_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n146)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h376C318CEC8017FF)) n147_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n147)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n148_lut (
        .I0(n144), .I1(n145), .I2(n146), .I3(n147), .I4(x[7]), .I5(x[10]), .O(n148)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n149_lut (
        .I0(n133), .I1(n138), .I2(n143), .I3(n148), .I4(x[3]), .I5(x[6]), .O(n149)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3D1F0A814F0A807E)) n150_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[9]), .O(n150)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3C033FF834BDFE81)) n151_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[9]), .O(n151)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5554338FCCC3C700)) n152_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[9]), .O(n152)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8002CCC32CE36300)) n153_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[8]), .I5(x[9]), .O(n153)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n154_lut (
        .I0(n150), .I1(n151), .I2(n152), .I3(n153), .I4(x[1]), .I5(x[10]), .O(n154)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n155_lut (
        .I0(~(n113)), .I1(~(n114)), .I2(~(n115)), .I3(~(n116)), .I4(x[1]), .I5(x[9]), .O(n155)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n156_lut (
        .I0(~(n118)), .I1(~(n119)), .I2(~(n120)), .I3(~(n121)), .I4(x[4]), .I5(x[9]), .O(n156)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n157_lut (
        .I0(~(n123)), .I1(~(n124)), .I2(~(n125)), .I3(~(n126)), .I4(x[1]), .I5(x[9]), .O(n157)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n158_lut (
        .I0(n154), .I1(n155), .I2(n156), .I3(n157), .I4(x[3]), .I5(x[7]), .O(n158)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n159_lut (
        .I0(~(n129)), .I1(~(n130)), .I2(~(n131)), .I3(~(n132)), .I4(x[8]), .I5(x[10]), .O(n159)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n160_lut (
        .I0(~(n134)), .I1(~(n135)), .I2(~(n136)), .I3(~(n137)), .I4(x[4]), .I5(x[8]), .O(n160)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n161_lut (
        .I0(~(n139)), .I1(~(n140)), .I2(~(n141)), .I3(~(n142)), .I4(x[4]), .I5(x[10]), .O(n161)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n162_lut (
        .I0(~(n144)), .I1(~(n145)), .I2(~(n146)), .I3(~(n147)), .I4(x[7]), .I5(x[10]), .O(n162)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n163_lut (
        .I0(n159), .I1(n160), .I2(n161), .I3(n162), .I4(x[3]), .I5(x[6]), .O(n163)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n164_lut (
        .I0(n128), .I1(n149), .I2(n158), .I3(n163), .I4(x[2]), .I5(x[11]), .O(n164)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE03FFC3E1F3EF0C0)) n165_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n165)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h013F03F01F1F7CF8)) n166_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n166)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h80F0FFF0F8FFFFFF)) n167_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n167)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8000FF00000000FF)) n168_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n168)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n169_lut (
        .I0(n165), .I1(n166), .I2(n167), .I3(n168), .I4(x[6]), .I5(x[10]), .O(n169)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC0E0E0C0C183071F)) n170_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n170)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC007FC03F03F0781)) n171_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n171)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3FFF7F00F801FFFF)) n172_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n172)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC08000C0FC0FF000)) n173_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n173)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n174_lut (
        .I0(n170), .I1(n171), .I2(n172), .I3(n173), .I4(x[8]), .I5(x[10]), .O(n174)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC037FF0FCFEFCF0)) n175_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n175)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hE0FC1F810FFC07C0)) n176_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n176)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC18181C000000000)) n177_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n177)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7CF8F0C0FFFF00FF)) n178_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n178)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n179_lut (
        .I0(n175), .I1(n176), .I2(n177), .I3(n178), .I4(x[7]), .I5(x[8]), .O(n179)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF00FFFE0F00EE8)) n180_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n180)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF0FFFFF070FFFF)) n181_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n181)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h17FFEEEEFF18F0FC)) n182_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n182)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC0013373108F1E0F)) n183_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n183)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n184_lut (
        .I0(n180), .I1(n181), .I2(n182), .I3(n183), .I4(x[2]), .I5(x[10]), .O(n184)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n185_lut (
        .I0(n169), .I1(n174), .I2(n179), .I3(n184), .I4(x[4]), .I5(x[9]), .O(n185)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF3EC17C07)) n186_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n186)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF0000FF07F01FE0)) n187_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n187)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8C0010701030307)) n188_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n188)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8800F7F1F070301)) n189_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[10]), .O(n189)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n190_lut (
        .I0(n186), .I1(n187), .I2(n188), .I3(n189), .I4(x[6]), .I5(x[9]), .O(n190)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFF1FF8FCF8F8)) n191_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n191)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0001000007030307)) n192_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n192)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h03C0F81F001FE07F)) n193_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n193)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF87E1F811FFF00FE)) n194_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[6]), .I5(x[10]), .O(n194)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n195_lut (
        .I0(n191), .I1(n192), .I2(n193), .I3(n194), .I4(x[4]), .I5(x[9]), .O(n195)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F07FCFFFCF803F0)) n196_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n196)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0F0C0E03F01F00F)) n197_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n197)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h070F000100FF3FE0)) n198_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n198)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8F0077FFF01037E)) n199_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[6]), .I4(x[9]), .I5(x[10]), .O(n199)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n200_lut (
        .I0(n196), .I1(n197), .I2(n198), .I3(n199), .I4(x[4]), .I5(x[5]), .O(n200)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1F7FFCE0810F7EF0)) n201_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n201)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFF00003F)) n202_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n202)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1F3F7FFFFFFF7F1F)) n203_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n203)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h07F01FC03E837C07)) n204_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n204)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n205_lut (
        .I0(n201), .I1(n202), .I2(n203), .I3(n204), .I4(x[9]), .I5(x[10]), .O(n205)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n206_lut (
        .I0(n190), .I1(n195), .I2(n200), .I3(n205), .I4(x[7]), .I5(x[8]), .O(n206)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1FC003C1E0C10F3E)) n207_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[5]), .I4(x[7]), .I5(x[8]), .O(n207)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n208_lut (
        .I0(n207), .I1(~(n166)), .I2(~(n167)), .I3(~(n168)), .I4(x[6]), .I5(x[10]), .O(n208)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n209_lut (
        .I0(~(n170)), .I1(~(n171)), .I2(~(n172)), .I3(~(n173)), .I4(x[8]), .I5(x[10]), .O(n209)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n210_lut (
        .I0(~(n175)), .I1(~(n176)), .I2(~(n177)), .I3(~(n178)), .I4(x[7]), .I5(x[8]), .O(n210)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n211_lut (
        .I0(~(n180)), .I1(~(n181)), .I2(~(n182)), .I3(~(n183)), .I4(x[2]), .I5(x[10]), .O(n211)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n212_lut (
        .I0(n208), .I1(n209), .I2(n210), .I3(n211), .I4(x[4]), .I5(x[9]), .O(n212)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n213_lut (
        .I0(~(n186)), .I1(~(n187)), .I2(~(n188)), .I3(~(n189)), .I4(x[6]), .I5(x[9]), .O(n213)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n214_lut (
        .I0(~(n191)), .I1(~(n192)), .I2(~(n193)), .I3(~(n194)), .I4(x[4]), .I5(x[9]), .O(n214)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n215_lut (
        .I0(~(n196)), .I1(~(n197)), .I2(~(n198)), .I3(~(n199)), .I4(x[4]), .I5(x[5]), .O(n215)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n216_lut (
        .I0(~(n201)), .I1(~(n202)), .I2(~(n203)), .I3(~(n204)), .I4(x[9]), .I5(x[10]), .O(n216)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n217_lut (
        .I0(n213), .I1(n214), .I2(n215), .I3(n216), .I4(x[7]), .I5(x[8]), .O(n217)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n218_lut (
        .I0(n185), .I1(n206), .I2(n212), .I3(n217), .I4(x[3]), .I5(x[11]), .O(n218)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h30CFF01008003070)) n219_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n219)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF0FFFFF00F0F0F)) n220_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n220)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F03F0030F00FFFF)) n221_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n221)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0C0010100CCF70C3)) n222_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n222)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n223_lut (
        .I0(n219), .I1(n220), .I2(n221), .I3(n222), .I4(x[9]), .I5(x[10]), .O(n223)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFFCFCF8F0C)) n224_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n224)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0F0FC800FF00CCF)) n225_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n225)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hEFF00FF0F80FC1C3)) n226_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n226)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFCFCFCFFFF0FF1F)) n227_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n227)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n228_lut (
        .I0(n224), .I1(n225), .I2(n226), .I3(n227), .I4(x[8]), .I5(x[9]), .O(n228)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0FC3FFFF7F7EFCF)) n229_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n229)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F0FC03F0EF00CCF)) n230_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n230)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF7F00CF003FC0F0F)) n231_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n231)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF3F3EFEFFFFF0000)) n232_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[10]), .O(n232)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n233_lut (
        .I0(n229), .I1(n230), .I2(n231), .I3(n232), .I4(x[8]), .I5(x[9]), .O(n233)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8F1CCFF0303030F1)) n234_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n234)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00E0800F83E3)) n235_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n235)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0F0F00FFFFF0FFF)) n236_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n236)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0C103030300CCF30)) n237_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n237)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n238_lut (
        .I0(n234), .I1(n235), .I2(n236), .I3(n237), .I4(x[9]), .I5(x[10]), .O(n238)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n239_lut (
        .I0(n223), .I1(n228), .I2(n233), .I3(n238), .I4(x[3]), .I5(x[5]), .O(n239)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h1CF3300C0C0C0030)) n240_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n240)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8FC3F0030F00FFFF)) n241_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n241)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0E0C080C0FE730F3)) n242_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n242)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n243_lut (
        .I0(n240), .I1(n220), .I2(n241), .I3(n242), .I4(x[9]), .I5(x[10]), .O(n243)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF0F0FFFF01FFFE)) n244_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n244)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCC0F3CFF30FF0CC8)) n245_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n245)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3F300000FCC7F0FF)) n246_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n246)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFF7FF00FFF007FE)) n247_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[6]), .I3(x[8]), .I4(x[9]), .I5(x[10]), .O(n247)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n248_lut (
        .I0(n244), .I1(n245), .I2(n246), .I3(n247), .I4(x[4]), .I5(x[7]), .O(n248)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF03F1FFF0FEFF7EF)) n249_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n249)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC707F0FE0FF0F3F3)) n250_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n250)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF3F70FF000000F0F)) n251_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n251)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h30F3F370FFFF037E)) n252_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[8]), .I5(x[10]), .O(n252)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n253_lut (
        .I0(n249), .I1(n250), .I2(n251), .I3(n252), .I4(x[7]), .I5(x[9]), .O(n253)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hC70CF37010001030)) n254_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n254)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00F0C00FC1F0)) n255_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n255)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0C081030100EE71C)) n256_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n256)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n257_lut (
        .I0(n254), .I1(n255), .I2(n236), .I3(n256), .I4(x[9]), .I5(x[10]), .O(n257)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n258_lut (
        .I0(n243), .I1(n248), .I2(n253), .I3(n257), .I4(x[3]), .I5(x[5]), .O(n258)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hCF300FEFF7FFCF8E)) n259_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n259)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n260_lut (
        .I0(n259), .I1(~(n220)), .I2(~(n221)), .I3(~(n222)), .I4(x[9]), .I5(x[10]), .O(n260)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n261_lut (
        .I0(~(n224)), .I1(~(n225)), .I2(~(n226)), .I3(~(n227)), .I4(x[8]), .I5(x[9]), .O(n261)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n262_lut (
        .I0(~(n229)), .I1(~(n230)), .I2(~(n231)), .I3(~(n232)), .I4(x[8]), .I5(x[9]), .O(n262)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n263_lut (
        .I0(~(n234)), .I1(~(n235)), .I2(~(n236)), .I3(~(n237)), .I4(x[9]), .I5(x[10]), .O(n263)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n264_lut (
        .I0(n260), .I1(n261), .I2(n262), .I3(n263), .I4(x[3]), .I5(x[5]), .O(n264)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n265_lut (
        .I0(~(n240)), .I1(~(n220)), .I2(~(n241)), .I3(~(n242)), .I4(x[9]), .I5(x[10]), .O(n265)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n266_lut (
        .I0(~(n244)), .I1(~(n245)), .I2(~(n246)), .I3(~(n247)), .I4(x[4]), .I5(x[7]), .O(n266)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n267_lut (
        .I0(~(n249)), .I1(~(n250)), .I2(~(n251)), .I3(~(n252)), .I4(x[7]), .I5(x[9]), .O(n267)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n268_lut (
        .I0(~(n254)), .I1(~(n255)), .I2(~(n236)), .I3(~(n256)), .I4(x[9]), .I5(x[10]), .O(n268)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n269_lut (
        .I0(n265), .I1(n266), .I2(n267), .I3(n268), .I4(x[3]), .I5(x[5]), .O(n269)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n270_lut (
        .I0(n239), .I1(n258), .I2(n264), .I3(n269), .I4(x[1]), .I5(x[11]), .O(n270)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8000F80000000000)) n271_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n271)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF003F0000)) n272_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n272)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0000FFFFFFFF)) n273_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n273)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFC0FFC00000FFFF)) n274_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n274)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n275_lut (
        .I0(n271), .I1(n272), .I2(n273), .I3(n274), .I4(x[8]), .I5(x[10]), .O(n275)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8000FFFEFFFFFFE0)) n276_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n276)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF01FFFFFFFFFF)) n277_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n277)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFC01FFFFFFFFFFF)) n278_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n278)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h03FF0FFF0007FFFC)) n279_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n279)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n280_lut (
        .I0(n276), .I1(n277), .I2(n278), .I3(n279), .I4(x[9]), .I5(x[10]), .O(n280)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC00FFFFFFFFFFFF)) n281_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n281)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000FFFF)) n282_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n282)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h007FFF000000FE00)) n283_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n283)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00070003FFFF0000)) n284_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n284)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n285_lut (
        .I0(n281), .I1(n282), .I2(n283), .I3(n284), .I4(x[7]), .I5(x[9]), .O(n285)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFF0003)) n286_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n286)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFE00000000000000)) n287_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n287)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF000FFFFC000003F)) n288_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n288)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00FF80FFFFFFF8)) n289_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n289)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n290_lut (
        .I0(n286), .I1(n287), .I2(n288), .I3(n289), .I4(x[7]), .I5(x[8]), .O(n290)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n291_lut (
        .I0(n275), .I1(n280), .I2(n285), .I3(n290), .I4(x[4]), .I5(x[6]), .O(n291)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3FFFFFFF03FF01FF)) n292_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n292)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF8000007FFFF001F)) n293_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n293)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000000000FF)) n294_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n294)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8000FFFFFFFFFFFF)) n295_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[9]), .I5(x[10]), .O(n295)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n296_lut (
        .I0(n292), .I1(n293), .I2(n294), .I3(n295), .I4(x[7]), .I5(x[8]), .O(n296)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFF8000C000)) n297_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n297)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FF000001FFFC00)) n298_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n298)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFE000000000000)) n299_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n299)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFF007F)) n300_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[8]), .I5(x[10]), .O(n300)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n301_lut (
        .I0(n297), .I1(n298), .I2(n299), .I3(n300), .I4(x[7]), .I5(x[9]), .O(n301)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF0300FFF0FFE080)) n302_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n302)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00FFFFFF07FFFF)) n303_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n303)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFF00)) n304_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n304)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0FFFFFFFFFFF7FC0)) n305_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[7]), .I4(x[9]), .I5(x[10]), .O(n305)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n306_lut (
        .I0(n302), .I1(n303), .I2(n304), .I3(n305), .I4(x[3]), .I5(x[8]), .O(n306)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFF07FF07FF)) n307_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n307)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFF0000)) n308_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n308)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h003F0003FFFFFFFF)) n309_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n309)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000010000F800)) n310_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[8]), .O(n310)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n311_lut (
        .I0(n307), .I1(n308), .I2(n309), .I3(n310), .I4(x[9]), .I5(x[10]), .O(n311)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n312_lut (
        .I0(n296), .I1(n301), .I2(n306), .I3(n311), .I4(x[4]), .I5(x[6]), .O(n312)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFF07FFFFFFFFFE)) n313_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n313)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n314_lut (
        .I0(n313), .I1(~(n272)), .I2(~(n273)), .I3(~(n274)), .I4(x[8]), .I5(x[10]), .O(n314)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n315_lut (
        .I0(~(n276)), .I1(~(n277)), .I2(~(n278)), .I3(~(n279)), .I4(x[9]), .I5(x[10]), .O(n315)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n316_lut (
        .I0(~(n281)), .I1(~(n282)), .I2(~(n283)), .I3(~(n284)), .I4(x[7]), .I5(x[9]), .O(n316)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n317_lut (
        .I0(~(n286)), .I1(~(n287)), .I2(~(n288)), .I3(~(n289)), .I4(x[7]), .I5(x[8]), .O(n317)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n318_lut (
        .I0(n314), .I1(n315), .I2(n316), .I3(n317), .I4(x[4]), .I5(x[6]), .O(n318)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n319_lut (
        .I0(~(n292)), .I1(~(n293)), .I2(~(n294)), .I3(~(n295)), .I4(x[7]), .I5(x[8]), .O(n319)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n320_lut (
        .I0(~(n297)), .I1(~(n298)), .I2(~(n299)), .I3(~(n300)), .I4(x[7]), .I5(x[9]), .O(n320)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n321_lut (
        .I0(~(n302)), .I1(~(n303)), .I2(~(n304)), .I3(~(n305)), .I4(x[3]), .I5(x[8]), .O(n321)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n322_lut (
        .I0(~(n307)), .I1(~(n308)), .I2(~(n309)), .I3(~(n310)), .I4(x[9]), .I5(x[10]), .O(n322)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n323_lut (
        .I0(n319), .I1(n320), .I2(n321), .I3(n322), .I4(x[4]), .I5(x[6]), .O(n323)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n324_lut (
        .I0(n291), .I1(n312), .I2(n318), .I3(n323), .I4(x[5]), .I5(x[11]), .O(n324)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFFFE000000)) n325_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n325)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0000001FFFFF)) n326_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n326)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00FFFFFFFFFFFFFF)) n327_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n327)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n328_lut (
        .I0(n325), .I1(n326), .I2(1'b1), .I3(n327), .I4(x[7]), .I5(x[10]), .O(n328)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000FF000000)) n329_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n329)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFC000000FFFF)) n330_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n330)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFFFFFFFFC0)) n331_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n331)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF000080000000)) n332_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n332)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n333_lut (
        .I0(n329), .I1(n330), .I2(n331), .I3(n332), .I4(x[6]), .I5(x[7]), .O(n333)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF03FFFFFF)) n334_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n334)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000F8000000)) n335_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n335)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF80000000000FFFF)) n336_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n336)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFFFFFFFF00)) n337_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n337)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n338_lut (
        .I0(n334), .I1(n335), .I2(n336), .I3(n337), .I4(x[6]), .I5(x[10]), .O(n338)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFC0FFFF0000)) n339_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n339)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF003FFFFFFFFF)) n340_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n340)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00008000FFFFFFFF)) n341_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n341)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n342_lut (
        .I0(n339), .I1(1'b1), .I2(n340), .I3(n341), .I4(x[5]), .I5(x[7]), .O(n342)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n343_lut (
        .I0(n328), .I1(n333), .I2(n338), .I3(n342), .I4(x[8]), .I5(x[9]), .O(n343)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF00030000)) n344_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n344)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFF800FFFF)) n345_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n345)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFF07FF0000)) n346_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[10]), .O(n346)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n347_lut (
        .I0(n344), .I1(n345), .I2(1'b1), .I3(n346), .I4(x[5]), .I5(x[7]), .O(n347)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h01FFFFFFFFFF0000)) n348_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n348)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00000000003F)) n349_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n349)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000003F00000000)) n350_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n350)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFF80FFFFFFFF)) n351_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[7]), .O(n351)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n352_lut (
        .I0(n348), .I1(n349), .I2(n350), .I3(n351), .I4(x[6]), .I5(x[10]), .O(n352)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000030000FFFF)) n353_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n353)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h07FFFFFFFFFF0000)) n354_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n354)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0000007FFFFF)) n355_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n355)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000001FF00000000)) n356_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[10]), .O(n356)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n357_lut (
        .I0(n353), .I1(n354), .I2(n355), .I3(n356), .I4(x[6]), .I5(x[7]), .O(n357)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFE00)) n358_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n358)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFF0000001FFFF)) n359_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n359)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000FFFFFF0000)) n360_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n360)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n361_lut (
        .I0(n358), .I1(1'b1), .I2(n359), .I3(n360), .I4(x[7]), .I5(x[10]), .O(n361)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n362_lut (
        .I0(n347), .I1(n352), .I2(n357), .I3(n361), .I4(x[8]), .I5(x[9]), .O(n362)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF000001FFFFFE)) n363_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[5]), .I5(x[6]), .O(n363)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n364_lut (
        .I0(n363), .I1(~(n326)), .I2(1'b0), .I3(~(n327)), .I4(x[7]), .I5(x[10]), .O(n364)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n365_lut (
        .I0(~(n329)), .I1(~(n330)), .I2(~(n331)), .I3(~(n332)), .I4(x[6]), .I5(x[7]), .O(n365)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n366_lut (
        .I0(~(n334)), .I1(~(n335)), .I2(~(n336)), .I3(~(n337)), .I4(x[6]), .I5(x[10]), .O(n366)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n367_lut (
        .I0(~(n339)), .I1(1'b0), .I2(~(n340)), .I3(~(n341)), .I4(x[5]), .I5(x[7]), .O(n367)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n368_lut (
        .I0(n364), .I1(n365), .I2(n366), .I3(n367), .I4(x[8]), .I5(x[9]), .O(n368)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n369_lut (
        .I0(~(n344)), .I1(~(n345)), .I2(1'b0), .I3(~(n346)), .I4(x[5]), .I5(x[7]), .O(n369)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n370_lut (
        .I0(~(n348)), .I1(~(n349)), .I2(~(n350)), .I3(~(n351)), .I4(x[6]), .I5(x[10]), .O(n370)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n371_lut (
        .I0(~(n353)), .I1(~(n354)), .I2(~(n355)), .I3(~(n356)), .I4(x[6]), .I5(x[7]), .O(n371)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n372_lut (
        .I0(~(n358)), .I1(1'b0), .I2(~(n359)), .I3(~(n360)), .I4(x[7]), .I5(x[10]), .O(n372)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n373_lut (
        .I0(n369), .I1(n370), .I2(n371), .I3(n372), .I4(x[8]), .I5(x[9]), .O(n373)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n374_lut (
        .I0(n343), .I1(n362), .I2(n368), .I3(n373), .I4(x[4]), .I5(x[11]), .O(n374)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000FFFFFFFF0000)) n375_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n375)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000003FF001F0000)) n376_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n376)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF000000000000)) n377_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n377)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n378_lut (
        .I0(n375), .I1(n376), .I2(n377), .I3(~(n375)), .I4(x[5]), .I5(x[6]), .O(n378)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0000FFFFFFFF)) n379_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[7]), .O(n379)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00000000FFFF)) n380_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[7]), .O(n380)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n381_lut (
        .I0(n379), .I1(n380), .I2(1'b1), .I3(1'b1), .I4(x[5]), .I5(x[9]), .O(n381)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF8000000FFFFF)) n382_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n382)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFF000000FFFFF)) n383_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n383)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n384_lut (
        .I0(1'b1), .I1(1'b1), .I2(n382), .I3(n383), .I4(x[2]), .I5(x[9]), .O(n384)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF003F0000FFFF)) n385_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n385)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7FFF00000000FFFF)) n386_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n386)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000000003FF)) n387_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n387)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n388_lut (
        .I0(n385), .I1(n386), .I2(n387), .I3(n375), .I4(x[5]), .I5(x[6]), .O(n388)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n389_lut (
        .I0(n378), .I1(n381), .I2(n384), .I3(n388), .I4(x[8]), .I5(x[10]), .O(n389)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF80000000000000)) n390_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n390)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00000000FFFC)) n391_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n391)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF0000F800FFFF)) n392_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n392)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n393_lut (
        .I0(n375), .I1(n390), .I2(n391), .I3(n392), .I4(x[5]), .I5(x[6]), .O(n393)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFE0000007FFFF)) n394_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n394)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFF0000007FFFF)) n395_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n395)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n396_lut (
        .I0(n394), .I1(n395), .I2(1'b1), .I3(1'b1), .I4(x[0]), .I5(x[9]), .O(n396)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF0000FFFF)) n397_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[6]), .I5(x[7]), .O(n397)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n398_lut (
        .I0(1'b1), .I1(1'b1), .I2(n380), .I3(n397), .I4(x[5]), .I5(x[9]), .O(n398)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h000000000000FFFF)) n399_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n399)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000F000FF800000)) n400_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n400)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n401_lut (
        .I0(~(n375)), .I1(n399), .I2(n400), .I3(n375), .I4(x[5]), .I5(x[6]), .O(n401)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n402_lut (
        .I0(n393), .I1(n396), .I2(n398), .I3(n401), .I4(x[8]), .I5(x[10]), .O(n402)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFF00000000FFFE)) n403_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[7]), .I5(x[9]), .O(n403)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n404_lut (
        .I0(n403), .I1(~(n376)), .I2(~(n377)), .I3(n375), .I4(x[5]), .I5(x[6]), .O(n404)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n405_lut (
        .I0(~(n379)), .I1(~(n380)), .I2(1'b0), .I3(1'b0), .I4(x[5]), .I5(x[9]), .O(n405)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n406_lut (
        .I0(1'b0), .I1(1'b0), .I2(~(n382)), .I3(~(n383)), .I4(x[2]), .I5(x[9]), .O(n406)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n407_lut (
        .I0(~(n385)), .I1(~(n386)), .I2(~(n387)), .I3(~(n375)), .I4(x[5]), .I5(x[6]), .O(n407)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n408_lut (
        .I0(n404), .I1(n405), .I2(n406), .I3(n407), .I4(x[8]), .I5(x[10]), .O(n408)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n409_lut (
        .I0(~(n375)), .I1(~(n390)), .I2(~(n391)), .I3(~(n392)), .I4(x[5]), .I5(x[6]), .O(n409)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n410_lut (
        .I0(~(n394)), .I1(~(n395)), .I2(1'b0), .I3(1'b0), .I4(x[0]), .I5(x[9]), .O(n410)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n411_lut (
        .I0(1'b0), .I1(1'b0), .I2(~(n380)), .I3(~(n397)), .I4(x[5]), .I5(x[9]), .O(n411)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n412_lut (
        .I0(n375), .I1(~(n399)), .I2(~(n400)), .I3(~(n375)), .I4(x[5]), .I5(x[6]), .O(n412)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n413_lut (
        .I0(n409), .I1(n410), .I2(n411), .I3(n412), .I4(x[8]), .I5(x[10]), .O(n413)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n414_lut (
        .I0(n389), .I1(n402), .I2(n408), .I3(n413), .I4(x[4]), .I5(x[11]), .O(n414)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFF00000000)) n415_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n415)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h003FFFFFFFFFFFFF)) n416_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n416)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n417_lut (
        .I0(1'b0), .I1(n415), .I2(n416), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n417)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n418_lut (
        .I0(n415), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n418)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h007FFFFFFFFFFFFF)) n419_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n419)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n420_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(n419), .I4(x[7]), .I5(x[8]), .O(n420)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0FFFFFFFFFFFFFFF)) n421_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n421)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n422_lut (
        .I0(1'b0), .I1(n415), .I2(n421), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n422)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n423_lut (
        .I0(n417), .I1(n418), .I2(n420), .I3(n422), .I4(x[9]), .I5(x[10]), .O(n423)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFFE0)) n424_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n424)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n425_lut (
        .I0(1'b0), .I1(n424), .I2(~(n415)), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n425)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFC00)) n426_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n426)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n427_lut (
        .I0(n426), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n427)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n428_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(~(n415)), .I4(x[7]), .I5(x[8]), .O(n428)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFF800)) n429_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n429)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n430_lut (
        .I0(1'b0), .I1(n429), .I2(~(n415)), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n430)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n431_lut (
        .I0(n425), .I1(n427), .I2(n428), .I3(n430), .I4(x[9]), .I5(x[10]), .O(n431)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFFFE)) n432_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[6]), .O(n432)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n433_lut (
        .I0(n432), .I1(~(n415)), .I2(~(n416)), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n433)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n434_lut (
        .I0(~(n415)), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n434)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n435_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(~(n419)), .I4(x[7]), .I5(x[8]), .O(n435)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n436_lut (
        .I0(1'b1), .I1(~(n415)), .I2(~(n421)), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n436)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n437_lut (
        .I0(n433), .I1(n434), .I2(n435), .I3(n436), .I4(x[9]), .I5(x[10]), .O(n437)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n438_lut (
        .I0(1'b1), .I1(~(n424)), .I2(n415), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n438)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n439_lut (
        .I0(~(n426)), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n439)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n440_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(n415), .I4(x[7]), .I5(x[8]), .O(n440)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n441_lut (
        .I0(1'b1), .I1(~(n429)), .I2(n415), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n441)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n442_lut (
        .I0(n438), .I1(n439), .I2(n440), .I3(n441), .I4(x[9]), .I5(x[10]), .O(n442)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n443_lut (
        .I0(n423), .I1(n431), .I2(n437), .I3(n442), .I4(x[5]), .I5(x[11]), .O(n443)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFF80000000000)) n444_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n444)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n445_lut (
        .I0(1'b0), .I1(1'b0), .I2(n444), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n445)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n446_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n446)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000003FFFFF)) n447_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n447)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n448_lut (
        .I0(1'b1), .I1(n447), .I2(1'b0), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n448)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n449_lut (
        .I0(n445), .I1(n446), .I2(n446), .I3(n448), .I4(x[9]), .I5(x[10]), .O(n449)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h00000000001FFFFF)) n450_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n450)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n451_lut (
        .I0(1'b1), .I1(n450), .I2(1'b0), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n451)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n452_lut (
        .I0(n445), .I1(n446), .I2(n446), .I3(n451), .I4(x[9]), .I5(x[10]), .O(n452)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFFFFFFFFFFFFFFFE)) n453_lut (
        .I0(x[1]), .I1(x[2]), .I2(x[3]), .I3(x[4]), .I4(x[5]), .I5(x[6]), .O(n453)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n454_lut (
        .I0(n453), .I1(1'b1), .I2(~(n444)), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n454)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n455_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n455)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n456_lut (
        .I0(1'b0), .I1(~(n447)), .I2(1'b1), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n456)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n457_lut (
        .I0(n454), .I1(n455), .I2(n455), .I3(n456), .I4(x[9]), .I5(x[10]), .O(n457)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n458_lut (
        .I0(1'b1), .I1(1'b1), .I2(~(n444)), .I3(1'b0), .I4(x[7]), .I5(x[8]), .O(n458)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n459_lut (
        .I0(1'b0), .I1(~(n450)), .I2(1'b1), .I3(1'b1), .I4(x[7]), .I5(x[8]), .O(n459)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n460_lut (
        .I0(n458), .I1(n455), .I2(n455), .I3(n459), .I4(x[9]), .I5(x[10]), .O(n460)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n461_lut (
        .I0(n449), .I1(n452), .I2(n457), .I3(n460), .I4(x[0]), .I5(x[11]), .O(n461)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n462_lut (
        .I0(1'b1), .I1(1'b1), .I2(1'b1), .I3(1'b1), .I4(x[6]), .I5(x[7]), .O(n462)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n463_lut (
        .I0(n462), .I1(n462), .I2(n462), .I3(n462), .I4(x[8]), .I5(x[9]), .O(n463)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0000000000000001)) n464_lut (
        .I0(x[0]), .I1(x[1]), .I2(x[2]), .I3(x[3]), .I4(x[4]), .I5(x[5]), .O(n464)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n465_lut (
        .I0(n464), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[7]), .O(n465)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n466_lut (
        .I0(1'b0), .I1(1'b0), .I2(1'b0), .I3(1'b0), .I4(x[6]), .I5(x[7]), .O(n466)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n467_lut (
        .I0(n465), .I1(n466), .I2(n466), .I3(n466), .I4(x[8]), .I5(x[9]), .O(n467)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n468_lut (
        .I0(n466), .I1(n466), .I2(n466), .I3(n466), .I4(x[8]), .I5(x[9]), .O(n468)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n469_lut (
        .I0(n463), .I1(n463), .I2(n467), .I3(n468), .I4(x[10]), .I5(x[11]), .O(n469)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA9593F3149A5965A)) n470_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n470)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h5A5A000E262596DA)) n471_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n471)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8C693800869B5A96)) n472_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n472)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h79D9C67CE1636AD6)) n473_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n473)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n474_lut (
        .I0(n470), .I1(n471), .I2(n472), .I3(n473), .I4(x[4]), .I5(x[6]), .O(n474)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h2FE8426C5585D5A5)) n475_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n475)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3CFFFFD3F57EAA5A)) n476_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n476)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0F9B185F334A55AA)) n477_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n477)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFC393368994B6A6A)) n478_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n478)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n479_lut (
        .I0(n475), .I1(n476), .I2(n477), .I3(n478), .I4(x[4]), .I5(x[6]), .O(n479)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA96999FFE255FD8F)) n480_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n480)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA95B3380792A00CF)) n481_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n481)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h256A87F41CB51527)) n482_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n482)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h695AC7FDF1B5954C)) n483_lut (
        .I0(x[0]), .I1(x[3]), .I2(x[4]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n483)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n484_lut (
        .I0(n480), .I1(n481), .I2(n482), .I3(n483), .I4(x[2]), .I5(x[6]), .O(n484)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h99699E1565A5D63E)) n485_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n485)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h66A4986AB9292B69)) n486_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n486)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h662AA64501000C0C)) n487_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n487)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hB9D55D9A3EF00F3C)) n488_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[9]), .O(n488)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n489_lut (
        .I0(n485), .I1(n486), .I2(n487), .I3(n488), .I4(x[3]), .I5(x[8]), .O(n489)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n490_lut (
        .I0(n474), .I1(n479), .I2(n484), .I3(n489), .I4(x[7]), .I5(x[10]), .O(n490)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0003583950074500)) n491_lut (
        .I0(x[4]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n491)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h015026C94DB4BAE7)) n492_lut (
        .I0(x[4]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n492)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h8780D631B1B8457E)) n493_lut (
        .I0(x[4]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n493)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hA69529F5F5C7B881)) n494_lut (
        .I0(x[4]), .I1(x[5]), .I2(x[6]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n494)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n495_lut (
        .I0(n491), .I1(n492), .I2(n493), .I3(n494), .I4(x[0]), .I5(x[2]), .O(n495)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h0B295A9A929617D5)) n496_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n496)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF0290D6576A65AAB)) n497_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n497)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h7C3C96B9BBABEAFF)) n498_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n498)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h3C137E962645688D)) n499_lut (
        .I0(x[0]), .I1(x[4]), .I2(x[5]), .I3(x[6]), .I4(x[7]), .I5(x[8]), .O(n499)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n500_lut (
        .I0(n496), .I1(n497), .I2(n498), .I3(n499), .I4(x[2]), .I5(x[10]), .O(n500)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h59596E93076AD3FC)) n501_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n501)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h66A9394020690F0F)) n502_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n502)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h666A490ACCA978F0)) n503_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n503)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h56A5B978FF79613C)) n504_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[7]), .I4(x[8]), .I5(x[10]), .O(n504)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n505_lut (
        .I0(n501), .I1(n502), .I2(n503), .I3(n504), .I4(x[5]), .I5(x[6]), .O(n505)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h668A0A0331300001)) n506_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n506)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hF00CDD00A9965A59)) n507_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n507)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h4469B9811A00FBC3)) n508_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n508)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hAB9999BA5A5AAA5A)) n509_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[4]), .I3(x[5]), .I4(x[6]), .I5(x[7]), .O(n509)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n510_lut (
        .I0(n506), .I1(n507), .I2(n508), .I3(n509), .I4(x[8]), .I5(x[10]), .O(n510)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n511_lut (
        .I0(n495), .I1(n500), .I2(n505), .I3(n510), .I4(x[3]), .I5(x[9]), .O(n511)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'h56A6C0CEB65A69A4)) n512_lut (
        .I0(x[0]), .I1(x[2]), .I2(x[3]), .I3(x[5]), .I4(x[8]), .I5(x[9]), .O(n512)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n513_lut (
        .I0(n512), .I1(~(n471)), .I2(~(n472)), .I3(~(n473)), .I4(x[4]), .I5(x[6]), .O(n513)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n514_lut (
        .I0(~(n475)), .I1(~(n476)), .I2(~(n477)), .I3(~(n478)), .I4(x[4]), .I5(x[6]), .O(n514)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n515_lut (
        .I0(~(n480)), .I1(~(n481)), .I2(~(n482)), .I3(~(n483)), .I4(x[2]), .I5(x[6]), .O(n515)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n516_lut (
        .I0(~(n485)), .I1(~(n486)), .I2(~(n487)), .I3(~(n488)), .I4(x[3]), .I5(x[8]), .O(n516)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n517_lut (
        .I0(n513), .I1(n514), .I2(n515), .I3(n516), .I4(x[7]), .I5(x[10]), .O(n517)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n518_lut (
        .I0(~(n491)), .I1(~(n492)), .I2(~(n493)), .I3(~(n494)), .I4(x[0]), .I5(x[2]), .O(n518)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n519_lut (
        .I0(~(n496)), .I1(~(n497)), .I2(~(n498)), .I3(~(n499)), .I4(x[2]), .I5(x[10]), .O(n519)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n520_lut (
        .I0(~(n501)), .I1(~(n502)), .I2(~(n503)), .I3(~(n504)), .I4(x[5]), .I5(x[6]), .O(n520)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n521_lut (
        .I0(~(n506)), .I1(~(n507)), .I2(~(n508)), .I3(~(n509)), .I4(x[8]), .I5(x[10]), .O(n521)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n522_lut (
        .I0(n518), .I1(n519), .I2(n520), .I3(n521), .I4(x[3]), .I5(x[9]), .O(n522)
    );

    (* DONT_TOUCH = "TRUE" *) plut_lut6 #(.INIT(64'hFF00F0F0CCCCAAAA)) n523_lut (
        .I0(n490), .I1(n511), .I2(n517), .I3(n522), .I4(x[1]), .I5(x[11]), .O(n523)
    );

    wire [10:0] ldtc_tss;
    wire [0:0] ldtc_td;
    assign ldtc_tss[0] = n53;
    assign ldtc_tss[1] = n107;
    assign ldtc_tss[2] = n164;
    assign ldtc_tss[3] = n218;
    assign ldtc_tss[4] = n270;
    assign ldtc_tss[5] = n324;
    assign ldtc_tss[6] = n374;
    assign ldtc_tss[7] = n414;
    assign ldtc_tss[8] = n443;
    assign ldtc_tss[9] = n461;
    assign ldtc_tss[10] = n469;
    assign ldtc_td[0] = n523;
    wire [11:0] ldtc_tss_ext = { { 1{1'b0} }, ldtc_tss } << 1;
    wire [11:0] ldtc_td_ext  = { { 11{1'b0} }, ldtc_td  };
    assign f = ldtc_tss_ext + ldtc_td_ext;
endmodule
